library IEEE;
use IEEE.std_logic_1164.all;
use work.SmartPackage.ALL;
use IEEE.numeric_std.all;

entity wallace_multiplier is
  port (
    a : in std_logic_vector(16 - 1 downto 0);
    b : in std_logic_vector(16 - 1 downto 0);
    c : out std_logic_vector(31 - 1 downto 0)
  );
end wallace_multiplier;

architecture Behavioral of wallace_multiplier is

    component full_adder is
     Port ( A : in STD_LOGIC;
             B : in STD_LOGIC;
             Cin : in STD_LOGIC;
             S : out STD_LOGIC;
             Cout : out STD_LOGIC);
    end component;

    component half_adder is
     Port ( A : in STD_LOGIC;
             B : in STD_LOGIC;
             S : out STD_LOGIC;
             Cout : out STD_LOGIC);
    end component;

    component carry_bypass_adder is
        Port ( A : in std_logic_vector(31 downto 0);
               B : in std_logic_vector(31 downto 0);
               S : out std_logic_vector(31 downto 0));
    end component;

    type partial_products_type is array (0 to 16 - 1) of std_logic_vector(16 - 1 downto 0);
    signal partial_products : partial_products_type;
    signal carry_bypass_a : std_logic_vector(31 downto 0);
    signal carry_bypass_b : std_logic_vector(31 downto 0);
    signal c_temp : std_logic_vector(31 downto 0);

    signal sum_764919 : std_logic;
signal cout_28774 : std_logic;
signal sum_579357 : std_logic;
signal cout_427899 : std_logic;
signal sum_786346 : std_logic;
signal cout_283914 : std_logic;
signal sum_822997 : std_logic;
signal cout_99255 : std_logic;
signal sum_222769 : std_logic;
signal cout_338740 : std_logic;
signal sum_494390 : std_logic;
signal cout_410342 : std_logic;
signal sum_557777 : std_logic;
signal cout_59262 : std_logic;
signal sum_180360 : std_logic;
signal cout_749781 : std_logic;
signal sum_410070 : std_logic;
signal cout_500237 : std_logic;
signal sum_101974 : std_logic;
signal cout_464992 : std_logic;
signal sum_275289 : std_logic;
signal cout_136981 : std_logic;
signal sum_952380 : std_logic;
signal cout_483752 : std_logic;
signal sum_568823 : std_logic;
signal cout_207780 : std_logic;
signal sum_147282 : std_logic;
signal cout_154835 : std_logic;
signal sum_916752 : std_logic;
signal cout_120483 : std_logic;
signal sum_826038 : std_logic;
signal cout_684194 : std_logic;
signal sum_827835 : std_logic;
signal cout_888683 : std_logic;
signal sum_490093 : std_logic;
signal cout_150064 : std_logic;
signal sum_651957 : std_logic;
signal cout_915659 : std_logic;
signal sum_702057 : std_logic;
signal cout_163734 : std_logic;
signal sum_251906 : std_logic;
signal cout_582835 : std_logic;
signal sum_160385 : std_logic;
signal cout_676755 : std_logic;
signal sum_100163 : std_logic;
signal cout_399438 : std_logic;
signal sum_519488 : std_logic;
signal cout_685880 : std_logic;
signal sum_948289 : std_logic;
signal cout_817181 : std_logic;
signal sum_275645 : std_logic;
signal cout_641831 : std_logic;
signal sum_905994 : std_logic;
signal cout_195612 : std_logic;
signal sum_471894 : std_logic;
signal cout_154881 : std_logic;
signal sum_902838 : std_logic;
signal cout_967259 : std_logic;
signal sum_855631 : std_logic;
signal cout_142187 : std_logic;
signal sum_404576 : std_logic;
signal cout_44885 : std_logic;
signal sum_241085 : std_logic;
signal cout_126830 : std_logic;
signal sum_439172 : std_logic;
signal cout_894990 : std_logic;
signal sum_750546 : std_logic;
signal cout_705138 : std_logic;
signal sum_269897 : std_logic;
signal cout_171096 : std_logic;
signal sum_565287 : std_logic;
signal cout_386117 : std_logic;
signal sum_822705 : std_logic;
signal cout_541205 : std_logic;
signal sum_800994 : std_logic;
signal cout_155961 : std_logic;
signal sum_252022 : std_logic;
signal cout_400811 : std_logic;
signal sum_417837 : std_logic;
signal cout_69827 : std_logic;
signal sum_325554 : std_logic;
signal cout_522329 : std_logic;
signal sum_15795 : std_logic;
signal cout_916594 : std_logic;
signal sum_369959 : std_logic;
signal cout_211052 : std_logic;
signal sum_541213 : std_logic;
signal cout_188951 : std_logic;
signal sum_129821 : std_logic;
signal cout_313582 : std_logic;
signal sum_733215 : std_logic;
signal cout_172496 : std_logic;
signal sum_257876 : std_logic;
signal cout_341273 : std_logic;
signal sum_76159 : std_logic;
signal cout_441877 : std_logic;
signal sum_800492 : std_logic;
signal cout_317830 : std_logic;
signal sum_649019 : std_logic;
signal cout_666012 : std_logic;
signal sum_401927 : std_logic;
signal cout_313956 : std_logic;
signal sum_764313 : std_logic;
signal cout_960814 : std_logic;
signal sum_509616 : std_logic;
signal cout_648745 : std_logic;
signal sum_874798 : std_logic;
signal cout_520934 : std_logic;
signal sum_290727 : std_logic;
signal cout_754725 : std_logic;
signal sum_785996 : std_logic;
signal cout_443029 : std_logic;
signal sum_757551 : std_logic;
signal cout_298758 : std_logic;
signal sum_860209 : std_logic;
signal cout_796262 : std_logic;
signal sum_564747 : std_logic;
signal cout_512704 : std_logic;
signal sum_781768 : std_logic;
signal cout_327114 : std_logic;
signal sum_49632 : std_logic;
signal cout_284124 : std_logic;
signal sum_374914 : std_logic;
signal cout_148635 : std_logic;
signal sum_811223 : std_logic;
signal cout_993789 : std_logic;
signal sum_627231 : std_logic;
signal cout_521027 : std_logic;
signal sum_859045 : std_logic;
signal cout_469424 : std_logic;
signal sum_368893 : std_logic;
signal cout_33075 : std_logic;
signal sum_921660 : std_logic;
signal cout_234614 : std_logic;
signal sum_395834 : std_logic;
signal cout_701326 : std_logic;
signal sum_551282 : std_logic;
signal cout_898933 : std_logic;
signal sum_107070 : std_logic;
signal cout_286406 : std_logic;
signal sum_564956 : std_logic;
signal cout_406130 : std_logic;
signal sum_214719 : std_logic;
signal cout_899981 : std_logic;
signal sum_553435 : std_logic;
signal cout_785622 : std_logic;
signal sum_525479 : std_logic;
signal cout_493344 : std_logic;
signal sum_190835 : std_logic;
signal cout_448862 : std_logic;
signal sum_742506 : std_logic;
signal cout_251932 : std_logic;
signal sum_511628 : std_logic;
signal cout_981885 : std_logic;
signal sum_256571 : std_logic;
signal cout_205302 : std_logic;
signal sum_187446 : std_logic;
signal cout_844520 : std_logic;
signal sum_499329 : std_logic;
signal cout_176804 : std_logic;
signal sum_794891 : std_logic;
signal cout_897676 : std_logic;
signal sum_570333 : std_logic;
signal cout_285129 : std_logic;
signal sum_376088 : std_logic;
signal cout_39979 : std_logic;
signal sum_978749 : std_logic;
signal cout_47287 : std_logic;
signal sum_156394 : std_logic;
signal cout_675045 : std_logic;
signal sum_143813 : std_logic;
signal cout_810133 : std_logic;
signal sum_412959 : std_logic;
signal cout_50814 : std_logic;
signal sum_89833 : std_logic;
signal cout_231264 : std_logic;
signal sum_352034 : std_logic;
signal cout_315014 : std_logic;
signal sum_480280 : std_logic;
signal cout_500323 : std_logic;
signal sum_833361 : std_logic;
signal cout_544773 : std_logic;
signal sum_752565 : std_logic;
signal cout_170918 : std_logic;
signal sum_954377 : std_logic;
signal cout_158710 : std_logic;
signal sum_707744 : std_logic;
signal cout_230667 : std_logic;
signal sum_536542 : std_logic;
signal cout_329486 : std_logic;
signal sum_845023 : std_logic;
signal cout_235510 : std_logic;
signal sum_870991 : std_logic;
signal cout_401666 : std_logic;
signal sum_199023 : std_logic;
signal cout_975011 : std_logic;
signal sum_273737 : std_logic;
signal cout_880735 : std_logic;
signal sum_142534 : std_logic;
signal cout_944096 : std_logic;
signal sum_510328 : std_logic;
signal cout_336691 : std_logic;
signal sum_665235 : std_logic;
signal cout_127219 : std_logic;
signal sum_697024 : std_logic;
signal cout_419323 : std_logic;
signal sum_257633 : std_logic;
signal cout_608182 : std_logic;
signal sum_382537 : std_logic;
signal cout_931374 : std_logic;
signal sum_161514 : std_logic;
signal cout_795340 : std_logic;
signal sum_969087 : std_logic;
signal cout_982442 : std_logic;
signal sum_767736 : std_logic;
signal cout_50397 : std_logic;
signal sum_100799 : std_logic;
signal cout_625517 : std_logic;
signal sum_232005 : std_logic;
signal cout_223032 : std_logic;
signal sum_878060 : std_logic;
signal cout_197320 : std_logic;
signal sum_606466 : std_logic;
signal cout_472778 : std_logic;
signal sum_385433 : std_logic;
signal cout_970632 : std_logic;
signal sum_667356 : std_logic;
signal cout_506445 : std_logic;
signal sum_683796 : std_logic;
signal cout_481211 : std_logic;
signal sum_305784 : std_logic;
signal cout_406184 : std_logic;
signal sum_554692 : std_logic;
signal cout_919075 : std_logic;
signal sum_570703 : std_logic;
signal cout_44492 : std_logic;
signal sum_722924 : std_logic;
signal cout_311266 : std_logic;
signal sum_268220 : std_logic;
signal cout_761351 : std_logic;
signal sum_402106 : std_logic;
signal cout_749422 : std_logic;
signal sum_409516 : std_logic;
signal cout_653208 : std_logic;
signal sum_661692 : std_logic;
signal cout_847021 : std_logic;
signal sum_367460 : std_logic;
signal cout_115092 : std_logic;
signal sum_951 : std_logic;
signal cout_524269 : std_logic;
signal sum_967160 : std_logic;
signal cout_507602 : std_logic;
signal sum_744015 : std_logic;
signal cout_323206 : std_logic;
signal sum_980106 : std_logic;
signal cout_945582 : std_logic;
signal sum_274585 : std_logic;
signal cout_452684 : std_logic;
signal sum_717014 : std_logic;
signal cout_679088 : std_logic;
signal sum_460096 : std_logic;
signal cout_224362 : std_logic;
signal sum_165640 : std_logic;
signal cout_111646 : std_logic;
signal sum_163022 : std_logic;
signal cout_858884 : std_logic;
signal sum_792035 : std_logic;
signal cout_30071 : std_logic;
signal sum_901306 : std_logic;
signal cout_956596 : std_logic;
signal sum_660823 : std_logic;
signal cout_868331 : std_logic;
signal sum_437656 : std_logic;
signal cout_416827 : std_logic;
signal sum_905681 : std_logic;
signal cout_435623 : std_logic;
signal sum_444952 : std_logic;
signal cout_476037 : std_logic;
signal sum_20721 : std_logic;
signal cout_201999 : std_logic;
signal sum_527568 : std_logic;
signal cout_539630 : std_logic;
signal sum_365635 : std_logic;
signal cout_874704 : std_logic;
signal sum_883412 : std_logic;
signal cout_300892 : std_logic;
signal sum_908827 : std_logic;
signal cout_414317 : std_logic;
signal sum_277432 : std_logic;
signal cout_618582 : std_logic;
signal sum_667288 : std_logic;
signal cout_564699 : std_logic;
signal sum_396396 : std_logic;
signal cout_372191 : std_logic;
signal sum_803175 : std_logic;
signal cout_713924 : std_logic;
signal sum_967664 : std_logic;
signal cout_75700 : std_logic;
signal sum_961901 : std_logic;
signal cout_571477 : std_logic;
signal sum_720232 : std_logic;
signal cout_339414 : std_logic;
signal sum_365138 : std_logic;
signal cout_74211 : std_logic;
signal sum_180499 : std_logic;
signal cout_113020 : std_logic;
signal sum_394816 : std_logic;
signal cout_991140 : std_logic;
signal sum_662358 : std_logic;
signal cout_732214 : std_logic;
signal sum_95985 : std_logic;
signal cout_592503 : std_logic;
signal sum_62223 : std_logic;
signal cout_808038 : std_logic;
signal sum_674809 : std_logic;
signal cout_997110 : std_logic;
signal sum_939359 : std_logic;
signal cout_193614 : std_logic;
signal sum_567775 : std_logic;
signal cout_983299 : std_logic;
signal sum_695865 : std_logic;
signal cout_658697 : std_logic;
signal sum_106498 : std_logic;
signal cout_987075 : std_logic;
signal sum_50326 : std_logic;
signal cout_197156 : std_logic;
signal sum_457415 : std_logic;
signal cout_81837 : std_logic;
signal sum_880909 : std_logic;
signal cout_588360 : std_logic;
signal sum_258244 : std_logic;
signal cout_384428 : std_logic;
signal sum_758416 : std_logic;
signal cout_772593 : std_logic;
signal sum_256046 : std_logic;
signal cout_956623 : std_logic;
signal sum_155656 : std_logic;
signal cout_968953 : std_logic;
signal sum_382851 : std_logic;
signal cout_213118 : std_logic;
signal sum_776758 : std_logic;
signal cout_31382 : std_logic;
signal sum_678538 : std_logic;
signal cout_720436 : std_logic;
signal sum_349666 : std_logic;
signal cout_186137 : std_logic;
signal sum_611747 : std_logic;
signal cout_775100 : std_logic;
signal sum_180812 : std_logic;
signal cout_605688 : std_logic;
signal sum_74962 : std_logic;
signal cout_806943 : std_logic;
signal sum_176515 : std_logic;
signal cout_688210 : std_logic;
signal sum_867437 : std_logic;
signal cout_660691 : std_logic;
signal sum_195682 : std_logic;
signal cout_55564 : std_logic;
signal sum_69528 : std_logic;
signal cout_284066 : std_logic;
signal sum_765424 : std_logic;
signal cout_550658 : std_logic;
signal sum_859277 : std_logic;
signal cout_12805 : std_logic;
signal sum_794561 : std_logic;
signal cout_616889 : std_logic;
signal sum_471696 : std_logic;
signal cout_966620 : std_logic;
signal sum_384372 : std_logic;
signal cout_50809 : std_logic;
signal sum_708540 : std_logic;
signal cout_136861 : std_logic;
signal sum_202319 : std_logic;
signal cout_438510 : std_logic;
signal sum_502356 : std_logic;
signal cout_698660 : std_logic;
signal sum_969478 : std_logic;
signal cout_78618 : std_logic;
signal sum_15498 : std_logic;
signal cout_332499 : std_logic;
signal sum_920500 : std_logic;
signal cout_639175 : std_logic;
signal sum_520498 : std_logic;
signal cout_411149 : std_logic;
signal sum_883481 : std_logic;
signal cout_341450 : std_logic;
signal sum_955207 : std_logic;
signal cout_347660 : std_logic;
signal sum_819480 : std_logic;
signal cout_862277 : std_logic;
signal sum_426993 : std_logic;
signal cout_585748 : std_logic;
signal sum_382685 : std_logic;
signal cout_985479 : std_logic;
signal sum_583731 : std_logic;
signal cout_365140 : std_logic;
signal sum_977460 : std_logic;
signal cout_861521 : std_logic;
signal sum_994015 : std_logic;
signal cout_551875 : std_logic;
signal sum_121008 : std_logic;
signal cout_406989 : std_logic;
signal sum_985669 : std_logic;
signal cout_358057 : std_logic;
signal sum_220091 : std_logic;
signal cout_826636 : std_logic;
signal sum_20111 : std_logic;
signal cout_579801 : std_logic;
signal sum_910987 : std_logic;
signal cout_185054 : std_logic;
signal sum_252974 : std_logic;
signal cout_688254 : std_logic;
signal sum_845494 : std_logic;
signal cout_682281 : std_logic;
signal sum_281821 : std_logic;
signal cout_837710 : std_logic;
signal sum_612520 : std_logic;
signal cout_43885 : std_logic;
signal sum_583673 : std_logic;
signal cout_609753 : std_logic;
signal pp_0_0 : std_logic;
signal pp_1_0 : std_logic;
signal pp_2_0 : std_logic;
signal pp_3_0 : std_logic;
signal pp_4_0 : std_logic;
signal pp_5_0 : std_logic;
signal pp_6_0 : std_logic;
signal pp_7_0 : std_logic;
signal pp_8_0 : std_logic;
signal pp_9_0 : std_logic;
signal pp_10_0 : std_logic;
signal pp_11_0 : std_logic;
signal pp_12_0 : std_logic;
signal pp_13_0 : std_logic;
signal pp_14_0 : std_logic;
signal pp_15_0 : std_logic;
signal pp_0_1 : std_logic;
signal pp_1_1 : std_logic;
signal pp_2_1 : std_logic;
signal pp_3_1 : std_logic;
signal pp_4_1 : std_logic;
signal pp_5_1 : std_logic;
signal pp_6_1 : std_logic;
signal pp_7_1 : std_logic;
signal pp_8_1 : std_logic;
signal pp_9_1 : std_logic;
signal pp_10_1 : std_logic;
signal pp_11_1 : std_logic;
signal pp_12_1 : std_logic;
signal pp_13_1 : std_logic;
signal pp_14_1 : std_logic;
signal pp_15_1 : std_logic;
signal pp_0_2 : std_logic;
signal pp_1_2 : std_logic;
signal pp_2_2 : std_logic;
signal pp_3_2 : std_logic;
signal pp_4_2 : std_logic;
signal pp_5_2 : std_logic;
signal pp_6_2 : std_logic;
signal pp_7_2 : std_logic;
signal pp_8_2 : std_logic;
signal pp_9_2 : std_logic;
signal pp_10_2 : std_logic;
signal pp_11_2 : std_logic;
signal pp_12_2 : std_logic;
signal pp_13_2 : std_logic;
signal pp_14_2 : std_logic;
signal pp_15_2 : std_logic;
signal pp_0_3 : std_logic;
signal pp_1_3 : std_logic;
signal pp_2_3 : std_logic;
signal pp_3_3 : std_logic;
signal pp_4_3 : std_logic;
signal pp_5_3 : std_logic;
signal pp_6_3 : std_logic;
signal pp_7_3 : std_logic;
signal pp_8_3 : std_logic;
signal pp_9_3 : std_logic;
signal pp_10_3 : std_logic;
signal pp_11_3 : std_logic;
signal pp_12_3 : std_logic;
signal pp_13_3 : std_logic;
signal pp_14_3 : std_logic;
signal pp_15_3 : std_logic;
signal pp_0_4 : std_logic;
signal pp_1_4 : std_logic;
signal pp_2_4 : std_logic;
signal pp_3_4 : std_logic;
signal pp_4_4 : std_logic;
signal pp_5_4 : std_logic;
signal pp_6_4 : std_logic;
signal pp_7_4 : std_logic;
signal pp_8_4 : std_logic;
signal pp_9_4 : std_logic;
signal pp_10_4 : std_logic;
signal pp_11_4 : std_logic;
signal pp_12_4 : std_logic;
signal pp_13_4 : std_logic;
signal pp_14_4 : std_logic;
signal pp_15_4 : std_logic;
signal pp_0_5 : std_logic;
signal pp_1_5 : std_logic;
signal pp_2_5 : std_logic;
signal pp_3_5 : std_logic;
signal pp_4_5 : std_logic;
signal pp_5_5 : std_logic;
signal pp_6_5 : std_logic;
signal pp_7_5 : std_logic;
signal pp_8_5 : std_logic;
signal pp_9_5 : std_logic;
signal pp_10_5 : std_logic;
signal pp_11_5 : std_logic;
signal pp_12_5 : std_logic;
signal pp_13_5 : std_logic;
signal pp_14_5 : std_logic;
signal pp_15_5 : std_logic;
signal pp_0_6 : std_logic;
signal pp_1_6 : std_logic;
signal pp_2_6 : std_logic;
signal pp_3_6 : std_logic;
signal pp_4_6 : std_logic;
signal pp_5_6 : std_logic;
signal pp_6_6 : std_logic;
signal pp_7_6 : std_logic;
signal pp_8_6 : std_logic;
signal pp_9_6 : std_logic;
signal pp_10_6 : std_logic;
signal pp_11_6 : std_logic;
signal pp_12_6 : std_logic;
signal pp_13_6 : std_logic;
signal pp_14_6 : std_logic;
signal pp_15_6 : std_logic;
signal pp_0_7 : std_logic;
signal pp_1_7 : std_logic;
signal pp_2_7 : std_logic;
signal pp_3_7 : std_logic;
signal pp_4_7 : std_logic;
signal pp_5_7 : std_logic;
signal pp_6_7 : std_logic;
signal pp_7_7 : std_logic;
signal pp_8_7 : std_logic;
signal pp_9_7 : std_logic;
signal pp_10_7 : std_logic;
signal pp_11_7 : std_logic;
signal pp_12_7 : std_logic;
signal pp_13_7 : std_logic;
signal pp_14_7 : std_logic;
signal pp_15_7 : std_logic;
signal pp_0_8 : std_logic;
signal pp_1_8 : std_logic;
signal pp_2_8 : std_logic;
signal pp_3_8 : std_logic;
signal pp_4_8 : std_logic;
signal pp_5_8 : std_logic;
signal pp_6_8 : std_logic;
signal pp_7_8 : std_logic;
signal pp_8_8 : std_logic;
signal pp_9_8 : std_logic;
signal pp_10_8 : std_logic;
signal pp_11_8 : std_logic;
signal pp_12_8 : std_logic;
signal pp_13_8 : std_logic;
signal pp_14_8 : std_logic;
signal pp_15_8 : std_logic;
signal pp_0_9 : std_logic;
signal pp_1_9 : std_logic;
signal pp_2_9 : std_logic;
signal pp_3_9 : std_logic;
signal pp_4_9 : std_logic;
signal pp_5_9 : std_logic;
signal pp_6_9 : std_logic;
signal pp_7_9 : std_logic;
signal pp_8_9 : std_logic;
signal pp_9_9 : std_logic;
signal pp_10_9 : std_logic;
signal pp_11_9 : std_logic;
signal pp_12_9 : std_logic;
signal pp_13_9 : std_logic;
signal pp_14_9 : std_logic;
signal pp_15_9 : std_logic;
signal pp_0_10 : std_logic;
signal pp_1_10 : std_logic;
signal pp_2_10 : std_logic;
signal pp_3_10 : std_logic;
signal pp_4_10 : std_logic;
signal pp_5_10 : std_logic;
signal pp_6_10 : std_logic;
signal pp_7_10 : std_logic;
signal pp_8_10 : std_logic;
signal pp_9_10 : std_logic;
signal pp_10_10 : std_logic;
signal pp_11_10 : std_logic;
signal pp_12_10 : std_logic;
signal pp_13_10 : std_logic;
signal pp_14_10 : std_logic;
signal pp_15_10 : std_logic;
signal pp_0_11 : std_logic;
signal pp_1_11 : std_logic;
signal pp_2_11 : std_logic;
signal pp_3_11 : std_logic;
signal pp_4_11 : std_logic;
signal pp_5_11 : std_logic;
signal pp_6_11 : std_logic;
signal pp_7_11 : std_logic;
signal pp_8_11 : std_logic;
signal pp_9_11 : std_logic;
signal pp_10_11 : std_logic;
signal pp_11_11 : std_logic;
signal pp_12_11 : std_logic;
signal pp_13_11 : std_logic;
signal pp_14_11 : std_logic;
signal pp_15_11 : std_logic;
signal pp_0_12 : std_logic;
signal pp_1_12 : std_logic;
signal pp_2_12 : std_logic;
signal pp_3_12 : std_logic;
signal pp_4_12 : std_logic;
signal pp_5_12 : std_logic;
signal pp_6_12 : std_logic;
signal pp_7_12 : std_logic;
signal pp_8_12 : std_logic;
signal pp_9_12 : std_logic;
signal pp_10_12 : std_logic;
signal pp_11_12 : std_logic;
signal pp_12_12 : std_logic;
signal pp_13_12 : std_logic;
signal pp_14_12 : std_logic;
signal pp_15_12 : std_logic;
signal pp_0_13 : std_logic;
signal pp_1_13 : std_logic;
signal pp_2_13 : std_logic;
signal pp_3_13 : std_logic;
signal pp_4_13 : std_logic;
signal pp_5_13 : std_logic;
signal pp_6_13 : std_logic;
signal pp_7_13 : std_logic;
signal pp_8_13 : std_logic;
signal pp_9_13 : std_logic;
signal pp_10_13 : std_logic;
signal pp_11_13 : std_logic;
signal pp_12_13 : std_logic;
signal pp_13_13 : std_logic;
signal pp_14_13 : std_logic;
signal pp_15_13 : std_logic;
signal pp_0_14 : std_logic;
signal pp_1_14 : std_logic;
signal pp_2_14 : std_logic;
signal pp_3_14 : std_logic;
signal pp_4_14 : std_logic;
signal pp_5_14 : std_logic;
signal pp_6_14 : std_logic;
signal pp_7_14 : std_logic;
signal pp_8_14 : std_logic;
signal pp_9_14 : std_logic;
signal pp_10_14 : std_logic;
signal pp_11_14 : std_logic;
signal pp_12_14 : std_logic;
signal pp_13_14 : std_logic;
signal pp_14_14 : std_logic;
signal pp_15_14 : std_logic;
signal pp_0_15 : std_logic;
signal pp_1_15 : std_logic;
signal pp_2_15 : std_logic;
signal pp_3_15 : std_logic;
signal pp_4_15 : std_logic;
signal pp_5_15 : std_logic;
signal pp_6_15 : std_logic;
signal pp_7_15 : std_logic;
signal pp_8_15 : std_logic;
signal pp_9_15 : std_logic;
signal pp_10_15 : std_logic;
signal pp_11_15 : std_logic;
signal pp_12_15 : std_logic;
signal pp_13_15 : std_logic;
signal pp_14_15 : std_logic;
signal pp_15_15 : std_logic;

begin

    c <= c_temp(30 downto 0);
    
        half_adder_36276 : half_adder
            port map (
                a => pp_0_15,
                b => pp_1_14,
                s => sum_764919,
                Cout => cout_28774
            );
        

        half_adder_38520 : half_adder
            port map (
                a => pp_1_15,
                b => pp_2_14,
                s => sum_579357,
                Cout => cout_427899
            );
        

        full_adder_66054 : full_adder
            port map (
                a => sum_764919,
                b => pp_2_13,
                Cin => pp_3_12,
                s => sum_822997,
                Cout => cout_99255
            );
        

        full_adder_91394 : full_adder
            port map (
                a => sum_579357,
                b => cout_28774,
                Cin => pp_3_13,
                s => sum_222769,
                Cout => cout_338740
            );
        

        full_adder_71145 : full_adder
            port map (
                a => cout_427899,
                b => pp_2_15,
                Cin => pp_3_14,
                s => sum_494390,
                Cout => cout_410342
            );
        

        half_adder_42921 : half_adder
            port map (
                a => pp_0_14,
                b => pp_1_13,
                s => sum_786346,
                Cout => cout_283914
            );
        

        full_adder_27921 : full_adder
            port map (
                a => sum_786346,
                b => pp_2_12,
                Cin => pp_3_11,
                s => sum_180360,
                Cout => cout_749781
            );
        

        full_adder_57093 : full_adder
            port map (
                a => sum_822997,
                b => cout_283914,
                Cin => pp_4_11,
                s => sum_410070,
                Cout => cout_500237
            );
        

        full_adder_30486 : full_adder
            port map (
                a => sum_222769,
                b => cout_99255,
                Cin => pp_4_12,
                s => sum_101974,
                Cout => cout_464992
            );
        

        full_adder_2654 : full_adder
            port map (
                a => sum_494390,
                b => cout_338740,
                Cin => pp_4_13,
                s => sum_275289,
                Cout => cout_136981
            );
        

        full_adder_26643 : full_adder
            port map (
                a => cout_410342,
                b => pp_3_15,
                Cin => pp_4_14,
                s => sum_952380,
                Cout => cout_483752
            );
        

        half_adder_80873 : half_adder
            port map (
                a => pp_0_13,
                b => pp_1_12,
                s => sum_557777,
                Cout => cout_59262
            );
        

        full_adder_95908 : full_adder
            port map (
                a => sum_557777,
                b => pp_2_11,
                Cin => pp_3_10,
                s => sum_147282,
                Cout => cout_154835
            );
        

        full_adder_85405 : full_adder
            port map (
                a => sum_180360,
                b => cout_59262,
                Cin => pp_4_10,
                s => sum_916752,
                Cout => cout_120483
            );
        

        full_adder_52860 : full_adder
            port map (
                a => sum_410070,
                b => cout_749781,
                Cin => pp_5_10,
                s => sum_826038,
                Cout => cout_684194
            );
        

        full_adder_94959 : full_adder
            port map (
                a => sum_101974,
                b => cout_500237,
                Cin => pp_5_11,
                s => sum_827835,
                Cout => cout_888683
            );
        

        full_adder_58855 : full_adder
            port map (
                a => sum_275289,
                b => cout_464992,
                Cin => pp_5_12,
                s => sum_490093,
                Cout => cout_150064
            );
        

        full_adder_21044 : full_adder
            port map (
                a => sum_952380,
                b => cout_136981,
                Cin => pp_5_13,
                s => sum_651957,
                Cout => cout_915659
            );
        

        full_adder_63133 : full_adder
            port map (
                a => cout_483752,
                b => pp_4_15,
                Cin => pp_5_14,
                s => sum_702057,
                Cout => cout_163734
            );
        

        half_adder_31535 : half_adder
            port map (
                a => pp_0_12,
                b => pp_1_11,
                s => sum_568823,
                Cout => cout_207780
            );
        

        full_adder_48321 : full_adder
            port map (
                a => sum_568823,
                b => pp_2_10,
                Cin => pp_3_9,
                s => sum_160385,
                Cout => cout_676755
            );
        

        full_adder_86208 : full_adder
            port map (
                a => sum_147282,
                b => cout_207780,
                Cin => pp_4_9,
                s => sum_100163,
                Cout => cout_399438
            );
        

        full_adder_28916 : full_adder
            port map (
                a => sum_916752,
                b => cout_154835,
                Cin => pp_5_9,
                s => sum_519488,
                Cout => cout_685880
            );
        

        full_adder_75163 : full_adder
            port map (
                a => sum_826038,
                b => cout_120483,
                Cin => pp_6_9,
                s => sum_948289,
                Cout => cout_817181
            );
        

        full_adder_61446 : full_adder
            port map (
                a => sum_827835,
                b => cout_684194,
                Cin => pp_6_10,
                s => sum_275645,
                Cout => cout_641831
            );
        

        full_adder_75364 : full_adder
            port map (
                a => sum_490093,
                b => cout_888683,
                Cin => pp_6_11,
                s => sum_905994,
                Cout => cout_195612
            );
        

        full_adder_391 : full_adder
            port map (
                a => sum_651957,
                b => cout_150064,
                Cin => pp_6_12,
                s => sum_471894,
                Cout => cout_154881
            );
        

        full_adder_48402 : full_adder
            port map (
                a => sum_702057,
                b => cout_915659,
                Cin => pp_6_13,
                s => sum_902838,
                Cout => cout_967259
            );
        

        full_adder_4376 : full_adder
            port map (
                a => cout_163734,
                b => pp_5_15,
                Cin => pp_6_14,
                s => sum_855631,
                Cout => cout_142187
            );
        

        half_adder_37221 : half_adder
            port map (
                a => pp_0_11,
                b => pp_1_10,
                s => sum_251906,
                Cout => cout_582835
            );
        

        full_adder_30369 : full_adder
            port map (
                a => sum_251906,
                b => pp_2_9,
                Cin => pp_3_8,
                s => sum_241085,
                Cout => cout_126830
            );
        

        full_adder_73504 : full_adder
            port map (
                a => sum_160385,
                b => cout_582835,
                Cin => pp_4_8,
                s => sum_439172,
                Cout => cout_894990
            );
        

        full_adder_95001 : full_adder
            port map (
                a => sum_100163,
                b => cout_676755,
                Cin => pp_5_8,
                s => sum_750546,
                Cout => cout_705138
            );
        

        full_adder_21951 : full_adder
            port map (
                a => sum_519488,
                b => cout_399438,
                Cin => pp_6_8,
                s => sum_269897,
                Cout => cout_171096
            );
        

        full_adder_37993 : full_adder
            port map (
                a => sum_948289,
                b => cout_685880,
                Cin => pp_7_8,
                s => sum_565287,
                Cout => cout_386117
            );
        

        full_adder_80758 : full_adder
            port map (
                a => sum_275645,
                b => cout_817181,
                Cin => pp_7_9,
                s => sum_822705,
                Cout => cout_541205
            );
        

        full_adder_71727 : full_adder
            port map (
                a => sum_905994,
                b => cout_641831,
                Cin => pp_7_10,
                s => sum_800994,
                Cout => cout_155961
            );
        

        full_adder_65250 : full_adder
            port map (
                a => sum_471894,
                b => cout_195612,
                Cin => pp_7_11,
                s => sum_252022,
                Cout => cout_400811
            );
        

        full_adder_40729 : full_adder
            port map (
                a => sum_902838,
                b => cout_154881,
                Cin => pp_7_12,
                s => sum_417837,
                Cout => cout_69827
            );
        

        full_adder_46493 : full_adder
            port map (
                a => sum_855631,
                b => cout_967259,
                Cin => pp_7_13,
                s => sum_325554,
                Cout => cout_522329
            );
        

        full_adder_61687 : full_adder
            port map (
                a => cout_142187,
                b => pp_6_15,
                Cin => pp_7_14,
                s => sum_15795,
                Cout => cout_916594
            );
        

        half_adder_3099 : half_adder
            port map (
                a => pp_0_10,
                b => pp_1_9,
                s => sum_404576,
                Cout => cout_44885
            );
        

        full_adder_99084 : full_adder
            port map (
                a => sum_404576,
                b => pp_2_8,
                Cin => pp_3_7,
                s => sum_541213,
                Cout => cout_188951
            );
        

        full_adder_8509 : full_adder
            port map (
                a => sum_241085,
                b => cout_44885,
                Cin => pp_4_7,
                s => sum_129821,
                Cout => cout_313582
            );
        

        full_adder_42648 : full_adder
            port map (
                a => sum_439172,
                b => cout_126830,
                Cin => pp_5_7,
                s => sum_733215,
                Cout => cout_172496
            );
        

        full_adder_93277 : full_adder
            port map (
                a => sum_750546,
                b => cout_894990,
                Cin => pp_6_7,
                s => sum_257876,
                Cout => cout_341273
            );
        

        full_adder_60704 : full_adder
            port map (
                a => sum_269897,
                b => cout_705138,
                Cin => pp_7_7,
                s => sum_76159,
                Cout => cout_441877
            );
        

        full_adder_16118 : full_adder
            port map (
                a => sum_565287,
                b => cout_171096,
                Cin => pp_8_7,
                s => sum_800492,
                Cout => cout_317830
            );
        

        full_adder_61289 : full_adder
            port map (
                a => sum_822705,
                b => cout_386117,
                Cin => pp_8_8,
                s => sum_649019,
                Cout => cout_666012
            );
        

        full_adder_22249 : full_adder
            port map (
                a => sum_800994,
                b => cout_541205,
                Cin => pp_8_9,
                s => sum_401927,
                Cout => cout_313956
            );
        

        full_adder_64740 : full_adder
            port map (
                a => sum_252022,
                b => cout_155961,
                Cin => pp_8_10,
                s => sum_764313,
                Cout => cout_960814
            );
        

        full_adder_47909 : full_adder
            port map (
                a => sum_417837,
                b => cout_400811,
                Cin => pp_8_11,
                s => sum_509616,
                Cout => cout_648745
            );
        

        full_adder_69968 : full_adder
            port map (
                a => sum_325554,
                b => cout_69827,
                Cin => pp_8_12,
                s => sum_874798,
                Cout => cout_520934
            );
        

        full_adder_23959 : full_adder
            port map (
                a => sum_15795,
                b => cout_522329,
                Cin => pp_8_13,
                s => sum_290727,
                Cout => cout_754725
            );
        

        full_adder_9793 : full_adder
            port map (
                a => cout_916594,
                b => pp_7_15,
                Cin => pp_8_14,
                s => sum_785996,
                Cout => cout_443029
            );
        

        half_adder_44099 : half_adder
            port map (
                a => pp_0_9,
                b => pp_1_8,
                s => sum_369959,
                Cout => cout_211052
            );
        

        full_adder_35112 : full_adder
            port map (
                a => sum_369959,
                b => pp_2_7,
                Cin => pp_3_6,
                s => sum_860209,
                Cout => cout_796262
            );
        

        full_adder_86692 : full_adder
            port map (
                a => sum_541213,
                b => cout_211052,
                Cin => pp_4_6,
                s => sum_564747,
                Cout => cout_512704
            );
        

        full_adder_39703 : full_adder
            port map (
                a => sum_129821,
                b => cout_188951,
                Cin => pp_5_6,
                s => sum_781768,
                Cout => cout_327114
            );
        

        full_adder_41857 : full_adder
            port map (
                a => sum_733215,
                b => cout_313582,
                Cin => pp_6_6,
                s => sum_49632,
                Cout => cout_284124
            );
        

        full_adder_15776 : full_adder
            port map (
                a => sum_257876,
                b => cout_172496,
                Cin => pp_7_6,
                s => sum_374914,
                Cout => cout_148635
            );
        

        full_adder_63622 : full_adder
            port map (
                a => sum_76159,
                b => cout_341273,
                Cin => pp_8_6,
                s => sum_811223,
                Cout => cout_993789
            );
        

        full_adder_92942 : full_adder
            port map (
                a => sum_800492,
                b => cout_441877,
                Cin => pp_9_6,
                s => sum_627231,
                Cout => cout_521027
            );
        

        full_adder_92987 : full_adder
            port map (
                a => sum_649019,
                b => cout_317830,
                Cin => pp_9_7,
                s => sum_859045,
                Cout => cout_469424
            );
        

        full_adder_59564 : full_adder
            port map (
                a => sum_401927,
                b => cout_666012,
                Cin => pp_9_8,
                s => sum_368893,
                Cout => cout_33075
            );
        

        full_adder_22651 : full_adder
            port map (
                a => sum_764313,
                b => cout_313956,
                Cin => pp_9_9,
                s => sum_921660,
                Cout => cout_234614
            );
        

        full_adder_91168 : full_adder
            port map (
                a => sum_509616,
                b => cout_960814,
                Cin => pp_9_10,
                s => sum_395834,
                Cout => cout_701326
            );
        

        full_adder_84775 : full_adder
            port map (
                a => sum_874798,
                b => cout_648745,
                Cin => pp_9_11,
                s => sum_551282,
                Cout => cout_898933
            );
        

        full_adder_75736 : full_adder
            port map (
                a => sum_290727,
                b => cout_520934,
                Cin => pp_9_12,
                s => sum_107070,
                Cout => cout_286406
            );
        

        full_adder_12319 : full_adder
            port map (
                a => sum_785996,
                b => cout_754725,
                Cin => pp_9_13,
                s => sum_564956,
                Cout => cout_406130
            );
        

        full_adder_19218 : full_adder
            port map (
                a => cout_443029,
                b => pp_8_15,
                Cin => pp_9_14,
                s => sum_214719,
                Cout => cout_899981
            );
        

        half_adder_82892 : half_adder
            port map (
                a => pp_0_8,
                b => pp_1_7,
                s => sum_757551,
                Cout => cout_298758
            );
        

        full_adder_15549 : full_adder
            port map (
                a => sum_757551,
                b => pp_2_6,
                Cin => pp_3_5,
                s => sum_525479,
                Cout => cout_493344
            );
        

        full_adder_69710 : full_adder
            port map (
                a => sum_860209,
                b => cout_298758,
                Cin => pp_4_5,
                s => sum_190835,
                Cout => cout_448862
            );
        

        full_adder_23759 : full_adder
            port map (
                a => sum_564747,
                b => cout_796262,
                Cin => pp_5_5,
                s => sum_742506,
                Cout => cout_251932
            );
        

        full_adder_89984 : full_adder
            port map (
                a => sum_781768,
                b => cout_512704,
                Cin => pp_6_5,
                s => sum_511628,
                Cout => cout_981885
            );
        

        full_adder_58454 : full_adder
            port map (
                a => sum_49632,
                b => cout_327114,
                Cin => pp_7_5,
                s => sum_256571,
                Cout => cout_205302
            );
        

        full_adder_73709 : full_adder
            port map (
                a => sum_374914,
                b => cout_284124,
                Cin => pp_8_5,
                s => sum_187446,
                Cout => cout_844520
            );
        

        full_adder_39197 : full_adder
            port map (
                a => sum_811223,
                b => cout_148635,
                Cin => pp_9_5,
                s => sum_499329,
                Cout => cout_176804
            );
        

        full_adder_59241 : full_adder
            port map (
                a => sum_627231,
                b => cout_993789,
                Cin => pp_10_5,
                s => sum_794891,
                Cout => cout_897676
            );
        

        full_adder_1163 : full_adder
            port map (
                a => sum_859045,
                b => cout_521027,
                Cin => pp_10_6,
                s => sum_570333,
                Cout => cout_285129
            );
        

        full_adder_8057 : full_adder
            port map (
                a => sum_368893,
                b => cout_469424,
                Cin => pp_10_7,
                s => sum_376088,
                Cout => cout_39979
            );
        

        full_adder_69950 : full_adder
            port map (
                a => sum_921660,
                b => cout_33075,
                Cin => pp_10_8,
                s => sum_978749,
                Cout => cout_47287
            );
        

        full_adder_88575 : full_adder
            port map (
                a => sum_395834,
                b => cout_234614,
                Cin => pp_10_9,
                s => sum_156394,
                Cout => cout_675045
            );
        

        full_adder_36450 : full_adder
            port map (
                a => sum_551282,
                b => cout_701326,
                Cin => pp_10_10,
                s => sum_143813,
                Cout => cout_810133
            );
        

        full_adder_87418 : full_adder
            port map (
                a => sum_107070,
                b => cout_898933,
                Cin => pp_10_11,
                s => sum_412959,
                Cout => cout_50814
            );
        

        full_adder_97047 : full_adder
            port map (
                a => sum_564956,
                b => cout_286406,
                Cin => pp_10_12,
                s => sum_89833,
                Cout => cout_231264
            );
        

        full_adder_47467 : full_adder
            port map (
                a => sum_214719,
                b => cout_406130,
                Cin => pp_10_13,
                s => sum_352034,
                Cout => cout_315014
            );
        

        full_adder_97869 : full_adder
            port map (
                a => cout_899981,
                b => pp_9_15,
                Cin => pp_10_14,
                s => sum_480280,
                Cout => cout_500323
            );
        

        half_adder_84238 : half_adder
            port map (
                a => pp_0_7,
                b => pp_1_6,
                s => sum_553435,
                Cout => cout_785622
            );
        

        full_adder_58988 : full_adder
            port map (
                a => sum_553435,
                b => pp_2_5,
                Cin => pp_3_4,
                s => sum_752565,
                Cout => cout_170918
            );
        

        full_adder_8967 : full_adder
            port map (
                a => sum_525479,
                b => cout_785622,
                Cin => pp_4_4,
                s => sum_954377,
                Cout => cout_158710
            );
        

        full_adder_33878 : full_adder
            port map (
                a => sum_190835,
                b => cout_493344,
                Cin => pp_5_4,
                s => sum_707744,
                Cout => cout_230667
            );
        

        full_adder_55907 : full_adder
            port map (
                a => sum_742506,
                b => cout_448862,
                Cin => pp_6_4,
                s => sum_536542,
                Cout => cout_329486
            );
        

        full_adder_23047 : full_adder
            port map (
                a => sum_511628,
                b => cout_251932,
                Cin => pp_7_4,
                s => sum_845023,
                Cout => cout_235510
            );
        

        full_adder_55015 : full_adder
            port map (
                a => sum_256571,
                b => cout_981885,
                Cin => pp_8_4,
                s => sum_870991,
                Cout => cout_401666
            );
        

        full_adder_75037 : full_adder
            port map (
                a => sum_187446,
                b => cout_205302,
                Cin => pp_9_4,
                s => sum_199023,
                Cout => cout_975011
            );
        

        full_adder_63052 : full_adder
            port map (
                a => sum_499329,
                b => cout_844520,
                Cin => pp_10_4,
                s => sum_273737,
                Cout => cout_880735
            );
        

        full_adder_2506 : full_adder
            port map (
                a => sum_794891,
                b => cout_176804,
                Cin => pp_11_4,
                s => sum_142534,
                Cout => cout_944096
            );
        

        full_adder_83292 : full_adder
            port map (
                a => sum_570333,
                b => cout_897676,
                Cin => pp_11_5,
                s => sum_510328,
                Cout => cout_336691
            );
        

        full_adder_32973 : full_adder
            port map (
                a => sum_376088,
                b => cout_285129,
                Cin => pp_11_6,
                s => sum_665235,
                Cout => cout_127219
            );
        

        full_adder_59130 : full_adder
            port map (
                a => sum_978749,
                b => cout_39979,
                Cin => pp_11_7,
                s => sum_697024,
                Cout => cout_419323
            );
        

        full_adder_83660 : full_adder
            port map (
                a => sum_156394,
                b => cout_47287,
                Cin => pp_11_8,
                s => sum_257633,
                Cout => cout_608182
            );
        

        full_adder_48538 : full_adder
            port map (
                a => sum_143813,
                b => cout_675045,
                Cin => pp_11_9,
                s => sum_382537,
                Cout => cout_931374
            );
        

        full_adder_88072 : full_adder
            port map (
                a => sum_412959,
                b => cout_810133,
                Cin => pp_11_10,
                s => sum_161514,
                Cout => cout_795340
            );
        

        full_adder_61452 : full_adder
            port map (
                a => sum_89833,
                b => cout_50814,
                Cin => pp_11_11,
                s => sum_969087,
                Cout => cout_982442
            );
        

        full_adder_31449 : full_adder
            port map (
                a => sum_352034,
                b => cout_231264,
                Cin => pp_11_12,
                s => sum_767736,
                Cout => cout_50397
            );
        

        full_adder_40572 : full_adder
            port map (
                a => sum_480280,
                b => cout_315014,
                Cin => pp_11_13,
                s => sum_100799,
                Cout => cout_625517
            );
        

        full_adder_64904 : full_adder
            port map (
                a => cout_500323,
                b => pp_10_15,
                Cin => pp_11_14,
                s => sum_232005,
                Cout => cout_223032
            );
        

        half_adder_89437 : half_adder
            port map (
                a => pp_0_6,
                b => pp_1_5,
                s => sum_833361,
                Cout => cout_544773
            );
        

        full_adder_63780 : full_adder
            port map (
                a => sum_833361,
                b => pp_2_4,
                Cin => pp_3_3,
                s => sum_606466,
                Cout => cout_472778
            );
        

        full_adder_31235 : full_adder
            port map (
                a => sum_752565,
                b => cout_544773,
                Cin => pp_4_3,
                s => sum_385433,
                Cout => cout_970632
            );
        

        full_adder_15929 : full_adder
            port map (
                a => sum_954377,
                b => cout_170918,
                Cin => pp_5_3,
                s => sum_667356,
                Cout => cout_506445
            );
        

        full_adder_38099 : full_adder
            port map (
                a => sum_707744,
                b => cout_158710,
                Cin => pp_6_3,
                s => sum_683796,
                Cout => cout_481211
            );
        

        full_adder_83466 : full_adder
            port map (
                a => sum_536542,
                b => cout_230667,
                Cin => pp_7_3,
                s => sum_305784,
                Cout => cout_406184
            );
        

        full_adder_6284 : full_adder
            port map (
                a => sum_845023,
                b => cout_329486,
                Cin => pp_8_3,
                s => sum_554692,
                Cout => cout_919075
            );
        

        full_adder_77952 : full_adder
            port map (
                a => sum_870991,
                b => cout_235510,
                Cin => pp_9_3,
                s => sum_570703,
                Cout => cout_44492
            );
        

        full_adder_98745 : full_adder
            port map (
                a => sum_199023,
                b => cout_401666,
                Cin => pp_10_3,
                s => sum_722924,
                Cout => cout_311266
            );
        

        full_adder_28122 : full_adder
            port map (
                a => sum_273737,
                b => cout_975011,
                Cin => pp_11_3,
                s => sum_268220,
                Cout => cout_761351
            );
        

        full_adder_23276 : full_adder
            port map (
                a => sum_142534,
                b => cout_880735,
                Cin => pp_12_3,
                s => sum_402106,
                Cout => cout_749422
            );
        

        full_adder_77508 : full_adder
            port map (
                a => sum_510328,
                b => cout_944096,
                Cin => pp_12_4,
                s => sum_409516,
                Cout => cout_653208
            );
        

        full_adder_63984 : full_adder
            port map (
                a => sum_665235,
                b => cout_336691,
                Cin => pp_12_5,
                s => sum_661692,
                Cout => cout_847021
            );
        

        full_adder_56462 : full_adder
            port map (
                a => sum_697024,
                b => cout_127219,
                Cin => pp_12_6,
                s => sum_367460,
                Cout => cout_115092
            );
        

        full_adder_57215 : full_adder
            port map (
                a => sum_257633,
                b => cout_419323,
                Cin => pp_12_7,
                s => sum_951,
                Cout => cout_524269
            );
        

        full_adder_514 : full_adder
            port map (
                a => sum_382537,
                b => cout_608182,
                Cin => pp_12_8,
                s => sum_967160,
                Cout => cout_507602
            );
        

        full_adder_58344 : full_adder
            port map (
                a => sum_161514,
                b => cout_931374,
                Cin => pp_12_9,
                s => sum_744015,
                Cout => cout_323206
            );
        

        full_adder_58923 : full_adder
            port map (
                a => sum_969087,
                b => cout_795340,
                Cin => pp_12_10,
                s => sum_980106,
                Cout => cout_945582
            );
        

        full_adder_65233 : full_adder
            port map (
                a => sum_767736,
                b => cout_982442,
                Cin => pp_12_11,
                s => sum_274585,
                Cout => cout_452684
            );
        

        full_adder_95442 : full_adder
            port map (
                a => sum_100799,
                b => cout_50397,
                Cin => pp_12_12,
                s => sum_717014,
                Cout => cout_679088
            );
        

        full_adder_31780 : full_adder
            port map (
                a => sum_232005,
                b => cout_625517,
                Cin => pp_12_13,
                s => sum_460096,
                Cout => cout_224362
            );
        

        full_adder_75609 : full_adder
            port map (
                a => cout_223032,
                b => pp_11_15,
                Cin => pp_12_14,
                s => sum_165640,
                Cout => cout_111646
            );
        

        half_adder_1895 : half_adder
            port map (
                a => pp_0_5,
                b => pp_1_4,
                s => sum_878060,
                Cout => cout_197320
            );
        

        full_adder_11925 : full_adder
            port map (
                a => sum_878060,
                b => pp_2_3,
                Cin => pp_3_2,
                s => sum_792035,
                Cout => cout_30071
            );
        

        full_adder_41844 : full_adder
            port map (
                a => sum_606466,
                b => cout_197320,
                Cin => pp_4_2,
                s => sum_901306,
                Cout => cout_956596
            );
        

        full_adder_29282 : full_adder
            port map (
                a => sum_385433,
                b => cout_472778,
                Cin => pp_5_2,
                s => sum_660823,
                Cout => cout_868331
            );
        

        full_adder_97547 : full_adder
            port map (
                a => sum_667356,
                b => cout_970632,
                Cin => pp_6_2,
                s => sum_437656,
                Cout => cout_416827
            );
        

        full_adder_50907 : full_adder
            port map (
                a => sum_683796,
                b => cout_506445,
                Cin => pp_7_2,
                s => sum_905681,
                Cout => cout_435623
            );
        

        full_adder_11618 : full_adder
            port map (
                a => sum_305784,
                b => cout_481211,
                Cin => pp_8_2,
                s => sum_444952,
                Cout => cout_476037
            );
        

        full_adder_65490 : full_adder
            port map (
                a => sum_554692,
                b => cout_406184,
                Cin => pp_9_2,
                s => sum_20721,
                Cout => cout_201999
            );
        

        full_adder_11336 : full_adder
            port map (
                a => sum_570703,
                b => cout_919075,
                Cin => pp_10_2,
                s => sum_527568,
                Cout => cout_539630
            );
        

        full_adder_77986 : full_adder
            port map (
                a => sum_722924,
                b => cout_44492,
                Cin => pp_11_2,
                s => sum_365635,
                Cout => cout_874704
            );
        

        full_adder_87421 : full_adder
            port map (
                a => sum_268220,
                b => cout_311266,
                Cin => pp_12_2,
                s => sum_883412,
                Cout => cout_300892
            );
        

        full_adder_62077 : full_adder
            port map (
                a => sum_402106,
                b => cout_761351,
                Cin => pp_13_2,
                s => sum_908827,
                Cout => cout_414317
            );
        

        full_adder_30936 : full_adder
            port map (
                a => sum_409516,
                b => cout_749422,
                Cin => pp_13_3,
                s => sum_277432,
                Cout => cout_618582
            );
        

        full_adder_14598 : full_adder
            port map (
                a => sum_661692,
                b => cout_653208,
                Cin => pp_13_4,
                s => sum_667288,
                Cout => cout_564699
            );
        

        full_adder_2053 : full_adder
            port map (
                a => sum_367460,
                b => cout_847021,
                Cin => pp_13_5,
                s => sum_396396,
                Cout => cout_372191
            );
        

        full_adder_22110 : full_adder
            port map (
                a => sum_951,
                b => cout_115092,
                Cin => pp_13_6,
                s => sum_803175,
                Cout => cout_713924
            );
        

        full_adder_3806 : full_adder
            port map (
                a => sum_967160,
                b => cout_524269,
                Cin => pp_13_7,
                s => sum_967664,
                Cout => cout_75700
            );
        

        full_adder_81165 : full_adder
            port map (
                a => sum_744015,
                b => cout_507602,
                Cin => pp_13_8,
                s => sum_961901,
                Cout => cout_571477
            );
        

        full_adder_60606 : full_adder
            port map (
                a => sum_980106,
                b => cout_323206,
                Cin => pp_13_9,
                s => sum_720232,
                Cout => cout_339414
            );
        

        full_adder_52276 : full_adder
            port map (
                a => sum_274585,
                b => cout_945582,
                Cin => pp_13_10,
                s => sum_365138,
                Cout => cout_74211
            );
        

        full_adder_64987 : full_adder
            port map (
                a => sum_717014,
                b => cout_452684,
                Cin => pp_13_11,
                s => sum_180499,
                Cout => cout_113020
            );
        

        full_adder_89593 : full_adder
            port map (
                a => sum_460096,
                b => cout_679088,
                Cin => pp_13_12,
                s => sum_394816,
                Cout => cout_991140
            );
        

        full_adder_88560 : full_adder
            port map (
                a => sum_165640,
                b => cout_224362,
                Cin => pp_13_13,
                s => sum_662358,
                Cout => cout_732214
            );
        

        full_adder_3692 : full_adder
            port map (
                a => cout_111646,
                b => pp_12_15,
                Cin => pp_13_14,
                s => sum_95985,
                Cout => cout_592503
            );
        

        half_adder_67530 : half_adder
            port map (
                a => pp_0_4,
                b => pp_1_3,
                s => sum_163022,
                Cout => cout_858884
            );
        

        full_adder_22118 : full_adder
            port map (
                a => sum_163022,
                b => pp_2_2,
                Cin => pp_3_1,
                s => sum_674809,
                Cout => cout_997110
            );
        

        full_adder_25601 : full_adder
            port map (
                a => sum_792035,
                b => cout_858884,
                Cin => pp_4_1,
                s => sum_939359,
                Cout => cout_193614
            );
        

        full_adder_49579 : full_adder
            port map (
                a => sum_901306,
                b => cout_30071,
                Cin => pp_5_1,
                s => sum_567775,
                Cout => cout_983299
            );
        

        full_adder_50338 : full_adder
            port map (
                a => sum_660823,
                b => cout_956596,
                Cin => pp_6_1,
                s => sum_695865,
                Cout => cout_658697
            );
        

        full_adder_313 : full_adder
            port map (
                a => sum_437656,
                b => cout_868331,
                Cin => pp_7_1,
                s => sum_106498,
                Cout => cout_987075
            );
        

        full_adder_94354 : full_adder
            port map (
                a => sum_905681,
                b => cout_416827,
                Cin => pp_8_1,
                s => sum_50326,
                Cout => cout_197156
            );
        

        full_adder_17070 : full_adder
            port map (
                a => sum_444952,
                b => cout_435623,
                Cin => pp_9_1,
                s => sum_457415,
                Cout => cout_81837
            );
        

        full_adder_49477 : full_adder
            port map (
                a => sum_20721,
                b => cout_476037,
                Cin => pp_10_1,
                s => sum_880909,
                Cout => cout_588360
            );
        

        full_adder_77334 : full_adder
            port map (
                a => sum_527568,
                b => cout_201999,
                Cin => pp_11_1,
                s => sum_258244,
                Cout => cout_384428
            );
        

        full_adder_23737 : full_adder
            port map (
                a => sum_365635,
                b => cout_539630,
                Cin => pp_12_1,
                s => sum_758416,
                Cout => cout_772593
            );
        

        full_adder_89074 : full_adder
            port map (
                a => sum_883412,
                b => cout_874704,
                Cin => pp_13_1,
                s => sum_256046,
                Cout => cout_956623
            );
        

        full_adder_62137 : full_adder
            port map (
                a => sum_908827,
                b => cout_300892,
                Cin => pp_14_1,
                s => sum_155656,
                Cout => cout_968953
            );
        

        full_adder_56430 : full_adder
            port map (
                a => sum_277432,
                b => cout_414317,
                Cin => pp_14_2,
                s => sum_382851,
                Cout => cout_213118
            );
        

        full_adder_66705 : full_adder
            port map (
                a => sum_667288,
                b => cout_618582,
                Cin => pp_14_3,
                s => sum_776758,
                Cout => cout_31382
            );
        

        full_adder_82420 : full_adder
            port map (
                a => sum_396396,
                b => cout_564699,
                Cin => pp_14_4,
                s => sum_678538,
                Cout => cout_720436
            );
        

        full_adder_77783 : full_adder
            port map (
                a => sum_803175,
                b => cout_372191,
                Cin => pp_14_5,
                s => sum_349666,
                Cout => cout_186137
            );
        

        full_adder_25259 : full_adder
            port map (
                a => sum_967664,
                b => cout_713924,
                Cin => pp_14_6,
                s => sum_611747,
                Cout => cout_775100
            );
        

        full_adder_7301 : full_adder
            port map (
                a => sum_961901,
                b => cout_75700,
                Cin => pp_14_7,
                s => sum_180812,
                Cout => cout_605688
            );
        

        full_adder_24544 : full_adder
            port map (
                a => sum_720232,
                b => cout_571477,
                Cin => pp_14_8,
                s => sum_74962,
                Cout => cout_806943
            );
        

        full_adder_70939 : full_adder
            port map (
                a => sum_365138,
                b => cout_339414,
                Cin => pp_14_9,
                s => sum_176515,
                Cout => cout_688210
            );
        

        full_adder_22095 : full_adder
            port map (
                a => sum_180499,
                b => cout_74211,
                Cin => pp_14_10,
                s => sum_867437,
                Cout => cout_660691
            );
        

        full_adder_47931 : full_adder
            port map (
                a => sum_394816,
                b => cout_113020,
                Cin => pp_14_11,
                s => sum_195682,
                Cout => cout_55564
            );
        

        full_adder_9874 : full_adder
            port map (
                a => sum_662358,
                b => cout_991140,
                Cin => pp_14_12,
                s => sum_69528,
                Cout => cout_284066
            );
        

        full_adder_72710 : full_adder
            port map (
                a => sum_95985,
                b => cout_732214,
                Cin => pp_14_13,
                s => sum_765424,
                Cout => cout_550658
            );
        

        full_adder_23597 : full_adder
            port map (
                a => cout_592503,
                b => pp_13_15,
                Cin => pp_14_14,
                s => sum_859277,
                Cout => cout_12805
            );
        

        half_adder_5515 : half_adder
            port map (
                a => pp_0_3,
                b => pp_1_2,
                s => sum_62223,
                Cout => cout_808038
            );
        

        full_adder_7765 : full_adder
            port map (
                a => sum_62223,
                b => pp_2_1,
                Cin => pp_3_0,
                s => sum_471696,
                Cout => cout_966620
            );
        

        full_adder_56641 : full_adder
            port map (
                a => sum_674809,
                b => cout_808038,
                Cin => pp_4_0,
                s => sum_384372,
                Cout => cout_50809
            );
        

        full_adder_76363 : full_adder
            port map (
                a => sum_939359,
                b => cout_997110,
                Cin => pp_5_0,
                s => sum_708540,
                Cout => cout_136861
            );
        

        full_adder_16469 : full_adder
            port map (
                a => sum_567775,
                b => cout_193614,
                Cin => pp_6_0,
                s => sum_202319,
                Cout => cout_438510
            );
        

        full_adder_46930 : full_adder
            port map (
                a => sum_695865,
                b => cout_983299,
                Cin => pp_7_0,
                s => sum_502356,
                Cout => cout_698660
            );
        

        full_adder_8342 : full_adder
            port map (
                a => sum_106498,
                b => cout_658697,
                Cin => pp_8_0,
                s => sum_969478,
                Cout => cout_78618
            );
        

        full_adder_21173 : full_adder
            port map (
                a => sum_50326,
                b => cout_987075,
                Cin => pp_9_0,
                s => sum_15498,
                Cout => cout_332499
            );
        

        full_adder_2162 : full_adder
            port map (
                a => sum_457415,
                b => cout_197156,
                Cin => pp_10_0,
                s => sum_920500,
                Cout => cout_639175
            );
        

        full_adder_87672 : full_adder
            port map (
                a => sum_880909,
                b => cout_81837,
                Cin => pp_11_0,
                s => sum_520498,
                Cout => cout_411149
            );
        

        full_adder_33396 : full_adder
            port map (
                a => sum_258244,
                b => cout_588360,
                Cin => pp_12_0,
                s => sum_883481,
                Cout => cout_341450
            );
        

        full_adder_39073 : full_adder
            port map (
                a => sum_758416,
                b => cout_384428,
                Cin => pp_13_0,
                s => sum_955207,
                Cout => cout_347660
            );
        

        full_adder_75719 : full_adder
            port map (
                a => sum_256046,
                b => cout_772593,
                Cin => pp_14_0,
                s => sum_819480,
                Cout => cout_862277
            );
        

        full_adder_80832 : full_adder
            port map (
                a => sum_155656,
                b => cout_956623,
                Cin => pp_15_0,
                s => sum_426993,
                Cout => cout_585748
            );
        

        full_adder_96319 : full_adder
            port map (
                a => sum_382851,
                b => cout_968953,
                Cin => pp_15_1,
                s => sum_382685,
                Cout => cout_985479
            );
        

        full_adder_2153 : full_adder
            port map (
                a => sum_776758,
                b => cout_213118,
                Cin => pp_15_2,
                s => sum_583731,
                Cout => cout_365140
            );
        

        full_adder_95539 : full_adder
            port map (
                a => sum_678538,
                b => cout_31382,
                Cin => pp_15_3,
                s => sum_977460,
                Cout => cout_861521
            );
        

        full_adder_5815 : full_adder
            port map (
                a => sum_349666,
                b => cout_720436,
                Cin => pp_15_4,
                s => sum_994015,
                Cout => cout_551875
            );
        

        full_adder_69159 : full_adder
            port map (
                a => sum_611747,
                b => cout_186137,
                Cin => pp_15_5,
                s => sum_121008,
                Cout => cout_406989
            );
        

        full_adder_19399 : full_adder
            port map (
                a => sum_180812,
                b => cout_775100,
                Cin => pp_15_6,
                s => sum_985669,
                Cout => cout_358057
            );
        

        full_adder_73786 : full_adder
            port map (
                a => sum_74962,
                b => cout_605688,
                Cin => pp_15_7,
                s => sum_220091,
                Cout => cout_826636
            );
        

        full_adder_97052 : full_adder
            port map (
                a => sum_176515,
                b => cout_806943,
                Cin => pp_15_8,
                s => sum_20111,
                Cout => cout_579801
            );
        

        full_adder_94460 : full_adder
            port map (
                a => sum_867437,
                b => cout_688210,
                Cin => pp_15_9,
                s => sum_910987,
                Cout => cout_185054
            );
        

        full_adder_30801 : full_adder
            port map (
                a => sum_195682,
                b => cout_660691,
                Cin => pp_15_10,
                s => sum_252974,
                Cout => cout_688254
            );
        

        full_adder_84307 : full_adder
            port map (
                a => sum_69528,
                b => cout_55564,
                Cin => pp_15_11,
                s => sum_845494,
                Cout => cout_682281
            );
        

        full_adder_86637 : full_adder
            port map (
                a => sum_765424,
                b => cout_284066,
                Cin => pp_15_12,
                s => sum_281821,
                Cout => cout_837710
            );
        

        full_adder_58853 : full_adder
            port map (
                a => sum_859277,
                b => cout_550658,
                Cin => pp_15_13,
                s => sum_612520,
                Cout => cout_43885
            );
        

        full_adder_51253 : full_adder
            port map (
                a => cout_12805,
                b => pp_14_15,
                Cin => pp_15_14,
                s => sum_583673,
                Cout => cout_609753
            );
        

        half_adder_58860 : half_adder
            port map (
                a => pp_0_2,
                b => pp_1_1,
                s => sum_794561,
                Cout => cout_616889
            );
        

        pp_0_0 <= a(0) and b(0);
        

        pp_1_0 <= a(1) and b(0);
        

        pp_2_0 <= a(2) and b(0);
        

        pp_3_0 <= a(3) and b(0);
        

        pp_4_0 <= a(4) and b(0);
        

        pp_5_0 <= a(5) and b(0);
        

        pp_6_0 <= a(6) and b(0);
        

        pp_7_0 <= a(7) and b(0);
        

        pp_8_0 <= a(8) and b(0);
        

        pp_9_0 <= a(9) and b(0);
        

        pp_10_0 <= a(10) and b(0);
        

        pp_11_0 <= a(11) and b(0);
        

        pp_12_0 <= a(12) and b(0);
        

        pp_13_0 <= a(13) and b(0);
        

        pp_14_0 <= a(14) and b(0);
        

        pp_15_0 <= a(15) and b(0);
        

        pp_0_1 <= a(0) and b(1);
        

        pp_1_1 <= a(1) and b(1);
        

        pp_2_1 <= a(2) and b(1);
        

        pp_3_1 <= a(3) and b(1);
        

        pp_4_1 <= a(4) and b(1);
        

        pp_5_1 <= a(5) and b(1);
        

        pp_6_1 <= a(6) and b(1);
        

        pp_7_1 <= a(7) and b(1);
        

        pp_8_1 <= a(8) and b(1);
        

        pp_9_1 <= a(9) and b(1);
        

        pp_10_1 <= a(10) and b(1);
        

        pp_11_1 <= a(11) and b(1);
        

        pp_12_1 <= a(12) and b(1);
        

        pp_13_1 <= a(13) and b(1);
        

        pp_14_1 <= a(14) and b(1);
        

        pp_15_1 <= a(15) and b(1);
        

        pp_0_2 <= a(0) and b(2);
        

        pp_1_2 <= a(1) and b(2);
        

        pp_2_2 <= a(2) and b(2);
        

        pp_3_2 <= a(3) and b(2);
        

        pp_4_2 <= a(4) and b(2);
        

        pp_5_2 <= a(5) and b(2);
        

        pp_6_2 <= a(6) and b(2);
        

        pp_7_2 <= a(7) and b(2);
        

        pp_8_2 <= a(8) and b(2);
        

        pp_9_2 <= a(9) and b(2);
        

        pp_10_2 <= a(10) and b(2);
        

        pp_11_2 <= a(11) and b(2);
        

        pp_12_2 <= a(12) and b(2);
        

        pp_13_2 <= a(13) and b(2);
        

        pp_14_2 <= a(14) and b(2);
        

        pp_15_2 <= a(15) and b(2);
        

        pp_0_3 <= a(0) and b(3);
        

        pp_1_3 <= a(1) and b(3);
        

        pp_2_3 <= a(2) and b(3);
        

        pp_3_3 <= a(3) and b(3);
        

        pp_4_3 <= a(4) and b(3);
        

        pp_5_3 <= a(5) and b(3);
        

        pp_6_3 <= a(6) and b(3);
        

        pp_7_3 <= a(7) and b(3);
        

        pp_8_3 <= a(8) and b(3);
        

        pp_9_3 <= a(9) and b(3);
        

        pp_10_3 <= a(10) and b(3);
        

        pp_11_3 <= a(11) and b(3);
        

        pp_12_3 <= a(12) and b(3);
        

        pp_13_3 <= a(13) and b(3);
        

        pp_14_3 <= a(14) and b(3);
        

        pp_15_3 <= a(15) and b(3);
        

        pp_0_4 <= a(0) and b(4);
        

        pp_1_4 <= a(1) and b(4);
        

        pp_2_4 <= a(2) and b(4);
        

        pp_3_4 <= a(3) and b(4);
        

        pp_4_4 <= a(4) and b(4);
        

        pp_5_4 <= a(5) and b(4);
        

        pp_6_4 <= a(6) and b(4);
        

        pp_7_4 <= a(7) and b(4);
        

        pp_8_4 <= a(8) and b(4);
        

        pp_9_4 <= a(9) and b(4);
        

        pp_10_4 <= a(10) and b(4);
        

        pp_11_4 <= a(11) and b(4);
        

        pp_12_4 <= a(12) and b(4);
        

        pp_13_4 <= a(13) and b(4);
        

        pp_14_4 <= a(14) and b(4);
        

        pp_15_4 <= a(15) and b(4);
        

        pp_0_5 <= a(0) and b(5);
        

        pp_1_5 <= a(1) and b(5);
        

        pp_2_5 <= a(2) and b(5);
        

        pp_3_5 <= a(3) and b(5);
        

        pp_4_5 <= a(4) and b(5);
        

        pp_5_5 <= a(5) and b(5);
        

        pp_6_5 <= a(6) and b(5);
        

        pp_7_5 <= a(7) and b(5);
        

        pp_8_5 <= a(8) and b(5);
        

        pp_9_5 <= a(9) and b(5);
        

        pp_10_5 <= a(10) and b(5);
        

        pp_11_5 <= a(11) and b(5);
        

        pp_12_5 <= a(12) and b(5);
        

        pp_13_5 <= a(13) and b(5);
        

        pp_14_5 <= a(14) and b(5);
        

        pp_15_5 <= a(15) and b(5);
        

        pp_0_6 <= a(0) and b(6);
        

        pp_1_6 <= a(1) and b(6);
        

        pp_2_6 <= a(2) and b(6);
        

        pp_3_6 <= a(3) and b(6);
        

        pp_4_6 <= a(4) and b(6);
        

        pp_5_6 <= a(5) and b(6);
        

        pp_6_6 <= a(6) and b(6);
        

        pp_7_6 <= a(7) and b(6);
        

        pp_8_6 <= a(8) and b(6);
        

        pp_9_6 <= a(9) and b(6);
        

        pp_10_6 <= a(10) and b(6);
        

        pp_11_6 <= a(11) and b(6);
        

        pp_12_6 <= a(12) and b(6);
        

        pp_13_6 <= a(13) and b(6);
        

        pp_14_6 <= a(14) and b(6);
        

        pp_15_6 <= a(15) and b(6);
        

        pp_0_7 <= a(0) and b(7);
        

        pp_1_7 <= a(1) and b(7);
        

        pp_2_7 <= a(2) and b(7);
        

        pp_3_7 <= a(3) and b(7);
        

        pp_4_7 <= a(4) and b(7);
        

        pp_5_7 <= a(5) and b(7);
        

        pp_6_7 <= a(6) and b(7);
        

        pp_7_7 <= a(7) and b(7);
        

        pp_8_7 <= a(8) and b(7);
        

        pp_9_7 <= a(9) and b(7);
        

        pp_10_7 <= a(10) and b(7);
        

        pp_11_7 <= a(11) and b(7);
        

        pp_12_7 <= a(12) and b(7);
        

        pp_13_7 <= a(13) and b(7);
        

        pp_14_7 <= a(14) and b(7);
        

        pp_15_7 <= a(15) and b(7);
        

        pp_0_8 <= a(0) and b(8);
        

        pp_1_8 <= a(1) and b(8);
        

        pp_2_8 <= a(2) and b(8);
        

        pp_3_8 <= a(3) and b(8);
        

        pp_4_8 <= a(4) and b(8);
        

        pp_5_8 <= a(5) and b(8);
        

        pp_6_8 <= a(6) and b(8);
        

        pp_7_8 <= a(7) and b(8);
        

        pp_8_8 <= a(8) and b(8);
        

        pp_9_8 <= a(9) and b(8);
        

        pp_10_8 <= a(10) and b(8);
        

        pp_11_8 <= a(11) and b(8);
        

        pp_12_8 <= a(12) and b(8);
        

        pp_13_8 <= a(13) and b(8);
        

        pp_14_8 <= a(14) and b(8);
        

        pp_15_8 <= a(15) and b(8);
        

        pp_0_9 <= a(0) and b(9);
        

        pp_1_9 <= a(1) and b(9);
        

        pp_2_9 <= a(2) and b(9);
        

        pp_3_9 <= a(3) and b(9);
        

        pp_4_9 <= a(4) and b(9);
        

        pp_5_9 <= a(5) and b(9);
        

        pp_6_9 <= a(6) and b(9);
        

        pp_7_9 <= a(7) and b(9);
        

        pp_8_9 <= a(8) and b(9);
        

        pp_9_9 <= a(9) and b(9);
        

        pp_10_9 <= a(10) and b(9);
        

        pp_11_9 <= a(11) and b(9);
        

        pp_12_9 <= a(12) and b(9);
        

        pp_13_9 <= a(13) and b(9);
        

        pp_14_9 <= a(14) and b(9);
        

        pp_15_9 <= a(15) and b(9);
        

        pp_0_10 <= a(0) and b(10);
        

        pp_1_10 <= a(1) and b(10);
        

        pp_2_10 <= a(2) and b(10);
        

        pp_3_10 <= a(3) and b(10);
        

        pp_4_10 <= a(4) and b(10);
        

        pp_5_10 <= a(5) and b(10);
        

        pp_6_10 <= a(6) and b(10);
        

        pp_7_10 <= a(7) and b(10);
        

        pp_8_10 <= a(8) and b(10);
        

        pp_9_10 <= a(9) and b(10);
        

        pp_10_10 <= a(10) and b(10);
        

        pp_11_10 <= a(11) and b(10);
        

        pp_12_10 <= a(12) and b(10);
        

        pp_13_10 <= a(13) and b(10);
        

        pp_14_10 <= a(14) and b(10);
        

        pp_15_10 <= a(15) and b(10);
        

        pp_0_11 <= a(0) and b(11);
        

        pp_1_11 <= a(1) and b(11);
        

        pp_2_11 <= a(2) and b(11);
        

        pp_3_11 <= a(3) and b(11);
        

        pp_4_11 <= a(4) and b(11);
        

        pp_5_11 <= a(5) and b(11);
        

        pp_6_11 <= a(6) and b(11);
        

        pp_7_11 <= a(7) and b(11);
        

        pp_8_11 <= a(8) and b(11);
        

        pp_9_11 <= a(9) and b(11);
        

        pp_10_11 <= a(10) and b(11);
        

        pp_11_11 <= a(11) and b(11);
        

        pp_12_11 <= a(12) and b(11);
        

        pp_13_11 <= a(13) and b(11);
        

        pp_14_11 <= a(14) and b(11);
        

        pp_15_11 <= a(15) and b(11);
        

        pp_0_12 <= a(0) and b(12);
        

        pp_1_12 <= a(1) and b(12);
        

        pp_2_12 <= a(2) and b(12);
        

        pp_3_12 <= a(3) and b(12);
        

        pp_4_12 <= a(4) and b(12);
        

        pp_5_12 <= a(5) and b(12);
        

        pp_6_12 <= a(6) and b(12);
        

        pp_7_12 <= a(7) and b(12);
        

        pp_8_12 <= a(8) and b(12);
        

        pp_9_12 <= a(9) and b(12);
        

        pp_10_12 <= a(10) and b(12);
        

        pp_11_12 <= a(11) and b(12);
        

        pp_12_12 <= a(12) and b(12);
        

        pp_13_12 <= a(13) and b(12);
        

        pp_14_12 <= a(14) and b(12);
        

        pp_15_12 <= a(15) and b(12);
        

        pp_0_13 <= a(0) and b(13);
        

        pp_1_13 <= a(1) and b(13);
        

        pp_2_13 <= a(2) and b(13);
        

        pp_3_13 <= a(3) and b(13);
        

        pp_4_13 <= a(4) and b(13);
        

        pp_5_13 <= a(5) and b(13);
        

        pp_6_13 <= a(6) and b(13);
        

        pp_7_13 <= a(7) and b(13);
        

        pp_8_13 <= a(8) and b(13);
        

        pp_9_13 <= a(9) and b(13);
        

        pp_10_13 <= a(10) and b(13);
        

        pp_11_13 <= a(11) and b(13);
        

        pp_12_13 <= a(12) and b(13);
        

        pp_13_13 <= a(13) and b(13);
        

        pp_14_13 <= a(14) and b(13);
        

        pp_15_13 <= a(15) and b(13);
        

        pp_0_14 <= a(0) and b(14);
        

        pp_1_14 <= a(1) and b(14);
        

        pp_2_14 <= a(2) and b(14);
        

        pp_3_14 <= a(3) and b(14);
        

        pp_4_14 <= a(4) and b(14);
        

        pp_5_14 <= a(5) and b(14);
        

        pp_6_14 <= a(6) and b(14);
        

        pp_7_14 <= a(7) and b(14);
        

        pp_8_14 <= a(8) and b(14);
        

        pp_9_14 <= a(9) and b(14);
        

        pp_10_14 <= a(10) and b(14);
        

        pp_11_14 <= a(11) and b(14);
        

        pp_12_14 <= a(12) and b(14);
        

        pp_13_14 <= a(13) and b(14);
        

        pp_14_14 <= a(14) and b(14);
        

        pp_15_14 <= a(15) and b(14);
        

        pp_0_15 <= a(0) and b(15);
        

        pp_1_15 <= a(1) and b(15);
        

        pp_2_15 <= a(2) and b(15);
        

        pp_3_15 <= a(3) and b(15);
        

        pp_4_15 <= a(4) and b(15);
        

        pp_5_15 <= a(5) and b(15);
        

        pp_6_15 <= a(6) and b(15);
        

        pp_7_15 <= a(7) and b(15);
        

        pp_8_15 <= a(8) and b(15);
        

        pp_9_15 <= a(9) and b(15);
        

        pp_10_15 <= a(10) and b(15);
        

        pp_11_15 <= a(11) and b(15);
        

        pp_12_15 <= a(12) and b(15);
        

        pp_13_15 <= a(13) and b(15);
        

        pp_14_15 <= a(14) and b(15);
        

        pp_15_15 <= a(15) and b(15);
        

        carry_bypass_adder_0 : carry_bypass_adder
            port map (
                a => carry_bypass_a,
                b => carry_bypass_b,
                s => c_temp
            );
        
carry_bypass_a <= '0' & pp_15_15 & cout_43885 & cout_837710 & cout_682281 & cout_688254 & cout_185054 & cout_579801 & cout_826636 & cout_358057 & cout_406989 & cout_551875 & cout_861521 & cout_365140 & cout_985479 & cout_585748 & cout_862277 & cout_347660 & cout_341450 & cout_411149 & cout_639175 & cout_332499 & cout_78618 & cout_698660 & cout_438510 & cout_136861 & cout_50809 & cout_966620 & cout_616889 & pp_2_0 & pp_1_0 & pp_0_0;
carry_bypass_b <= '0' & cout_609753 & sum_583673 & sum_612520 & sum_281821 & sum_845494 & sum_252974 & sum_910987 & sum_20111 & sum_220091 & sum_985669 & sum_121008 & sum_994015 & sum_977460 & sum_583731 & sum_382685 & sum_426993 & sum_819480 & sum_955207 & sum_883481 & sum_520498 & sum_920500 & sum_15498 & sum_969478 & sum_502356 & sum_202319 & sum_708540 & sum_384372 & sum_471696 & sum_794561 & pp_0_1 & '0';

end Behavioral;
