library IEEE;
use IEEE.std_logic_1164.all;

entity wallace_multiplier is
  port (
    a : in std_logic_vector(16 - 1 downto 0);
    b : in std_logic_vector(16 - 1 downto 0);
    c : out std_logic_vector(31 - 1 downto 0)
  );
end wallace_multiplier;

architecture Behavioral of wallace_multiplier is

    component full_adder is
     Port ( A : in STD_LOGIC;
             B : in STD_LOGIC;
             Cin : in STD_LOGIC;
             S : out STD_LOGIC;
             Cout : out STD_LOGIC);
    end component;

    component half_adder is
     Port ( A : in STD_LOGIC;
             B : in STD_LOGIC;
             S : out STD_LOGIC;
             Cout : out STD_LOGIC);
    end component;

    type partial_products_type is array (0 to 16 - 1) of std_logic_vector(16 - 1 downto 0);
    signal partial_products : partial_products_type;

    signal sum_757675 : std_logic;
signal cout_769389 : std_logic;
signal sum_932346 : std_logic;
signal cout_39739 : std_logic;
signal sum_754583 : std_logic;
signal cout_624584 : std_logic;
signal sum_659249 : std_logic;
signal cout_356642 : std_logic;
signal sum_47972 : std_logic;
signal cout_39813 : std_logic;
signal sum_753784 : std_logic;
signal cout_172689 : std_logic;
signal sum_560320 : std_logic;
signal cout_578344 : std_logic;
signal sum_538566 : std_logic;
signal cout_172686 : std_logic;
signal sum_756610 : std_logic;
signal cout_567486 : std_logic;
signal sum_914016 : std_logic;
signal cout_913439 : std_logic;
signal sum_13181 : std_logic;
signal cout_841917 : std_logic;
signal sum_977726 : std_logic;
signal cout_932234 : std_logic;
signal sum_910513 : std_logic;
signal cout_94920 : std_logic;
signal sum_226390 : std_logic;
signal cout_940010 : std_logic;
signal sum_766179 : std_logic;
signal cout_491530 : std_logic;
signal sum_146247 : std_logic;
signal cout_749783 : std_logic;
signal sum_722838 : std_logic;
signal cout_905765 : std_logic;
signal sum_86012 : std_logic;
signal cout_598245 : std_logic;
signal sum_492003 : std_logic;
signal cout_191038 : std_logic;
signal sum_618163 : std_logic;
signal cout_578246 : std_logic;
signal sum_123741 : std_logic;
signal cout_285703 : std_logic;
signal sum_990655 : std_logic;
signal cout_976970 : std_logic;
signal sum_671502 : std_logic;
signal cout_446076 : std_logic;
signal sum_411192 : std_logic;
signal cout_461391 : std_logic;
signal sum_249416 : std_logic;
signal cout_945951 : std_logic;
signal sum_686986 : std_logic;
signal cout_712188 : std_logic;
signal sum_277628 : std_logic;
signal cout_640546 : std_logic;
signal sum_287843 : std_logic;
signal cout_275866 : std_logic;
signal sum_625716 : std_logic;
signal cout_989486 : std_logic;
signal sum_375464 : std_logic;
signal cout_567696 : std_logic;
signal sum_327095 : std_logic;
signal cout_863399 : std_logic;
signal sum_222046 : std_logic;
signal cout_206738 : std_logic;
signal sum_7087 : std_logic;
signal cout_262915 : std_logic;
signal sum_413141 : std_logic;
signal cout_670764 : std_logic;
signal sum_380765 : std_logic;
signal cout_918132 : std_logic;
signal sum_913153 : std_logic;
signal cout_561087 : std_logic;
signal sum_390680 : std_logic;
signal cout_357374 : std_logic;
signal sum_616616 : std_logic;
signal cout_786530 : std_logic;
signal sum_863047 : std_logic;
signal cout_960948 : std_logic;
signal sum_774946 : std_logic;
signal cout_203266 : std_logic;
signal sum_961775 : std_logic;
signal cout_860843 : std_logic;
signal sum_451910 : std_logic;
signal cout_420673 : std_logic;
signal sum_208632 : std_logic;
signal cout_771281 : std_logic;
signal sum_274274 : std_logic;
signal cout_930231 : std_logic;
signal sum_194968 : std_logic;
signal cout_157897 : std_logic;
signal sum_24183 : std_logic;
signal cout_551891 : std_logic;
signal sum_349866 : std_logic;
signal cout_433248 : std_logic;
signal sum_797979 : std_logic;
signal cout_187818 : std_logic;
signal sum_427572 : std_logic;
signal cout_923055 : std_logic;
signal sum_797511 : std_logic;
signal cout_878210 : std_logic;
signal sum_409507 : std_logic;
signal cout_697098 : std_logic;
signal sum_181157 : std_logic;
signal cout_537561 : std_logic;
signal sum_315286 : std_logic;
signal cout_987740 : std_logic;
signal sum_404304 : std_logic;
signal cout_22433 : std_logic;
signal sum_383733 : std_logic;
signal cout_632990 : std_logic;
signal sum_360115 : std_logic;
signal cout_174525 : std_logic;
signal sum_230909 : std_logic;
signal cout_727671 : std_logic;
signal sum_372567 : std_logic;
signal cout_539978 : std_logic;
signal sum_246201 : std_logic;
signal cout_258710 : std_logic;
signal sum_903520 : std_logic;
signal cout_815001 : std_logic;
signal sum_774546 : std_logic;
signal cout_346012 : std_logic;
signal sum_960667 : std_logic;
signal cout_937613 : std_logic;
signal sum_705137 : std_logic;
signal cout_153737 : std_logic;
signal sum_149238 : std_logic;
signal cout_702253 : std_logic;
signal sum_388368 : std_logic;
signal cout_529839 : std_logic;
signal sum_419352 : std_logic;
signal cout_167953 : std_logic;
signal sum_796092 : std_logic;
signal cout_759053 : std_logic;
signal sum_135226 : std_logic;
signal cout_725574 : std_logic;
signal sum_165325 : std_logic;
signal cout_242304 : std_logic;
signal sum_669906 : std_logic;
signal cout_810450 : std_logic;
signal sum_711628 : std_logic;
signal cout_666929 : std_logic;
signal sum_410690 : std_logic;
signal cout_22372 : std_logic;
signal sum_310349 : std_logic;
signal cout_82769 : std_logic;
signal sum_905500 : std_logic;
signal cout_525986 : std_logic;
signal sum_975960 : std_logic;
signal cout_263090 : std_logic;
signal sum_21048 : std_logic;
signal cout_649712 : std_logic;
signal sum_592564 : std_logic;
signal cout_366028 : std_logic;
signal sum_272977 : std_logic;
signal cout_69885 : std_logic;
signal sum_387065 : std_logic;
signal cout_272868 : std_logic;
signal sum_182442 : std_logic;
signal cout_922087 : std_logic;
signal sum_409 : std_logic;
signal cout_821655 : std_logic;
signal sum_808671 : std_logic;
signal cout_61302 : std_logic;
signal sum_113860 : std_logic;
signal cout_327241 : std_logic;
signal sum_248889 : std_logic;
signal cout_82325 : std_logic;
signal sum_343072 : std_logic;
signal cout_791728 : std_logic;
signal sum_659836 : std_logic;
signal cout_684959 : std_logic;
signal sum_658736 : std_logic;
signal cout_846804 : std_logic;
signal sum_241703 : std_logic;
signal cout_974942 : std_logic;
signal sum_324032 : std_logic;
signal cout_889121 : std_logic;
signal sum_647575 : std_logic;
signal cout_904012 : std_logic;
signal sum_742414 : std_logic;
signal cout_276204 : std_logic;
signal sum_641583 : std_logic;
signal cout_199542 : std_logic;
signal sum_752893 : std_logic;
signal cout_936261 : std_logic;
signal sum_548921 : std_logic;
signal cout_138274 : std_logic;
signal sum_461182 : std_logic;
signal cout_599211 : std_logic;
signal sum_319630 : std_logic;
signal cout_152176 : std_logic;
signal sum_533069 : std_logic;
signal cout_111262 : std_logic;
signal sum_887964 : std_logic;
signal cout_284285 : std_logic;
signal sum_835449 : std_logic;
signal cout_139640 : std_logic;
signal sum_993754 : std_logic;
signal cout_177382 : std_logic;
signal sum_504281 : std_logic;
signal cout_5038 : std_logic;
signal sum_909922 : std_logic;
signal cout_662043 : std_logic;
signal sum_766402 : std_logic;
signal cout_63167 : std_logic;
signal sum_439931 : std_logic;
signal cout_599694 : std_logic;
signal sum_911256 : std_logic;
signal cout_952902 : std_logic;
signal sum_530689 : std_logic;
signal cout_606994 : std_logic;
signal sum_442354 : std_logic;
signal cout_738496 : std_logic;
signal sum_85078 : std_logic;
signal cout_43875 : std_logic;
signal sum_716697 : std_logic;
signal cout_180198 : std_logic;
signal sum_579393 : std_logic;
signal cout_401825 : std_logic;
signal sum_964352 : std_logic;
signal cout_5705 : std_logic;
signal sum_878840 : std_logic;
signal cout_413325 : std_logic;
signal sum_952338 : std_logic;
signal cout_227086 : std_logic;
signal sum_922115 : std_logic;
signal cout_232219 : std_logic;
signal sum_584013 : std_logic;
signal cout_403061 : std_logic;
signal sum_859480 : std_logic;
signal cout_928577 : std_logic;
signal sum_807794 : std_logic;
signal cout_847359 : std_logic;
signal sum_202927 : std_logic;
signal cout_299193 : std_logic;
signal sum_830004 : std_logic;
signal cout_599178 : std_logic;
signal sum_418595 : std_logic;
signal cout_717070 : std_logic;
signal sum_877555 : std_logic;
signal cout_186640 : std_logic;
signal sum_885640 : std_logic;
signal cout_744469 : std_logic;
signal sum_568950 : std_logic;
signal cout_217500 : std_logic;
signal sum_37576 : std_logic;
signal cout_543060 : std_logic;
signal sum_871425 : std_logic;
signal cout_380034 : std_logic;
signal sum_963006 : std_logic;
signal cout_960555 : std_logic;
signal sum_179806 : std_logic;
signal cout_909674 : std_logic;
signal sum_622556 : std_logic;
signal cout_6366 : std_logic;
signal sum_100853 : std_logic;
signal cout_241998 : std_logic;
signal sum_590812 : std_logic;
signal cout_189105 : std_logic;
signal sum_853972 : std_logic;
signal cout_908865 : std_logic;
signal sum_487151 : std_logic;
signal cout_428500 : std_logic;
signal sum_151833 : std_logic;
signal cout_442253 : std_logic;
signal sum_190083 : std_logic;
signal cout_44270 : std_logic;
signal sum_155461 : std_logic;
signal cout_752478 : std_logic;
signal sum_70271 : std_logic;
signal cout_103199 : std_logic;
signal sum_325561 : std_logic;
signal cout_503461 : std_logic;
signal sum_384618 : std_logic;
signal cout_554463 : std_logic;
signal sum_610884 : std_logic;
signal cout_963328 : std_logic;
signal sum_527017 : std_logic;
signal cout_836750 : std_logic;
signal sum_330037 : std_logic;
signal cout_845115 : std_logic;
signal sum_617507 : std_logic;
signal cout_187919 : std_logic;
signal sum_745173 : std_logic;
signal cout_903116 : std_logic;
signal sum_107552 : std_logic;
signal cout_57875 : std_logic;
signal sum_3669 : std_logic;
signal cout_924814 : std_logic;
signal sum_890133 : std_logic;
signal cout_752540 : std_logic;
signal sum_285660 : std_logic;
signal cout_750878 : std_logic;
signal sum_865435 : std_logic;
signal cout_347189 : std_logic;
signal sum_165169 : std_logic;
signal cout_903701 : std_logic;
signal sum_161296 : std_logic;
signal cout_9966 : std_logic;
signal sum_210485 : std_logic;
signal cout_154367 : std_logic;
signal sum_940061 : std_logic;
signal cout_777808 : std_logic;
signal sum_556282 : std_logic;
signal cout_918370 : std_logic;
signal sum_409267 : std_logic;
signal cout_765436 : std_logic;
signal sum_16716 : std_logic;
signal cout_743533 : std_logic;
signal sum_128628 : std_logic;
signal cout_809894 : std_logic;
signal sum_393354 : std_logic;
signal cout_773384 : std_logic;
signal sum_491221 : std_logic;
signal cout_681963 : std_logic;
signal sum_372577 : std_logic;
signal cout_12222 : std_logic;
signal sum_352335 : std_logic;
signal cout_194219 : std_logic;
signal sum_218632 : std_logic;
signal cout_283181 : std_logic;
signal sum_509457 : std_logic;
signal cout_801902 : std_logic;
signal sum_813250 : std_logic;
signal cout_597879 : std_logic;
signal sum_436895 : std_logic;
signal cout_52308 : std_logic;
signal sum_608641 : std_logic;
signal cout_230642 : std_logic;
signal sum_75594 : std_logic;
signal cout_269720 : std_logic;
signal sum_538112 : std_logic;
signal cout_612378 : std_logic;
signal sum_752554 : std_logic;
signal cout_390278 : std_logic;
signal sum_447835 : std_logic;
signal cout_81863 : std_logic;
signal sum_604064 : std_logic;
signal cout_665374 : std_logic;
signal sum_602802 : std_logic;
signal cout_313284 : std_logic;
signal sum_447776 : std_logic;
signal cout_610447 : std_logic;
signal sum_846479 : std_logic;
signal cout_58374 : std_logic;
signal sum_175238 : std_logic;
signal cout_352004 : std_logic;
signal sum_101042 : std_logic;
signal cout_120477 : std_logic;
signal sum_863612 : std_logic;
signal cout_621744 : std_logic;
signal sum_292728 : std_logic;
signal cout_253376 : std_logic;
signal sum_36423 : std_logic;
signal cout_986139 : std_logic;
signal sum_763057 : std_logic;
signal cout_830405 : std_logic;
signal sum_677725 : std_logic;
signal cout_225273 : std_logic;
signal sum_924856 : std_logic;
signal cout_105480 : std_logic;
signal sum_653807 : std_logic;
signal cout_683444 : std_logic;
signal sum_652062 : std_logic;
signal cout_734723 : std_logic;
signal sum_454017 : std_logic;
signal cout_648852 : std_logic;
signal sum_615388 : std_logic;
signal cout_622190 : std_logic;
signal sum_307052 : std_logic;
signal cout_296984 : std_logic;
signal sum_957721 : std_logic;
signal cout_372708 : std_logic;
signal sum_910907 : std_logic;
signal cout_87182 : std_logic;
signal sum_190554 : std_logic;
signal cout_901791 : std_logic;
signal sum_108552 : std_logic;
signal cout_938354 : std_logic;
signal sum_871398 : std_logic;
signal cout_899840 : std_logic;
signal sum_748543 : std_logic;
signal cout_473235 : std_logic;
signal sum_620884 : std_logic;
signal cout_502572 : std_logic;
signal sum_835826 : std_logic;
signal cout_615799 : std_logic;
signal sum_747437 : std_logic;
signal cout_907232 : std_logic;
signal sum_408519 : std_logic;
signal cout_273843 : std_logic;
signal sum_825709 : std_logic;
signal cout_593623 : std_logic;
signal sum_751602 : std_logic;
signal cout_860894 : std_logic;
signal sum_739794 : std_logic;
signal cout_336777 : std_logic;
signal sum_422751 : std_logic;
signal cout_174675 : std_logic;
signal sum_573526 : std_logic;
signal cout_622573 : std_logic;
signal sum_334672 : std_logic;
signal cout_614796 : std_logic;
signal sum_445479 : std_logic;
signal cout_694665 : std_logic;
signal sum_873056 : std_logic;
signal cout_34362 : std_logic;
signal sum_860833 : std_logic;
signal cout_288058 : std_logic;
signal sum_906512 : std_logic;
signal cout_430498 : std_logic;
signal sum_319921 : std_logic;
signal cout_310125 : std_logic;
signal sum_777791 : std_logic;
signal cout_278529 : std_logic;
signal sum_134521 : std_logic;
signal cout_907380 : std_logic;
signal sum_453295 : std_logic;
signal cout_505573 : std_logic;
signal pp_0_0 : std_logic;
signal pp_1_0 : std_logic;
signal pp_2_0 : std_logic;
signal pp_3_0 : std_logic;
signal pp_4_0 : std_logic;
signal pp_5_0 : std_logic;
signal pp_6_0 : std_logic;
signal pp_7_0 : std_logic;
signal pp_8_0 : std_logic;
signal pp_9_0 : std_logic;
signal pp_10_0 : std_logic;
signal pp_11_0 : std_logic;
signal pp_12_0 : std_logic;
signal pp_13_0 : std_logic;
signal pp_14_0 : std_logic;
signal pp_15_0 : std_logic;
signal pp_0_1 : std_logic;
signal pp_1_1 : std_logic;
signal pp_2_1 : std_logic;
signal pp_3_1 : std_logic;
signal pp_4_1 : std_logic;
signal pp_5_1 : std_logic;
signal pp_6_1 : std_logic;
signal pp_7_1 : std_logic;
signal pp_8_1 : std_logic;
signal pp_9_1 : std_logic;
signal pp_10_1 : std_logic;
signal pp_11_1 : std_logic;
signal pp_12_1 : std_logic;
signal pp_13_1 : std_logic;
signal pp_14_1 : std_logic;
signal pp_15_1 : std_logic;
signal pp_0_2 : std_logic;
signal pp_1_2 : std_logic;
signal pp_2_2 : std_logic;
signal pp_3_2 : std_logic;
signal pp_4_2 : std_logic;
signal pp_5_2 : std_logic;
signal pp_6_2 : std_logic;
signal pp_7_2 : std_logic;
signal pp_8_2 : std_logic;
signal pp_9_2 : std_logic;
signal pp_10_2 : std_logic;
signal pp_11_2 : std_logic;
signal pp_12_2 : std_logic;
signal pp_13_2 : std_logic;
signal pp_14_2 : std_logic;
signal pp_15_2 : std_logic;
signal pp_0_3 : std_logic;
signal pp_1_3 : std_logic;
signal pp_2_3 : std_logic;
signal pp_3_3 : std_logic;
signal pp_4_3 : std_logic;
signal pp_5_3 : std_logic;
signal pp_6_3 : std_logic;
signal pp_7_3 : std_logic;
signal pp_8_3 : std_logic;
signal pp_9_3 : std_logic;
signal pp_10_3 : std_logic;
signal pp_11_3 : std_logic;
signal pp_12_3 : std_logic;
signal pp_13_3 : std_logic;
signal pp_14_3 : std_logic;
signal pp_15_3 : std_logic;
signal pp_0_4 : std_logic;
signal pp_1_4 : std_logic;
signal pp_2_4 : std_logic;
signal pp_3_4 : std_logic;
signal pp_4_4 : std_logic;
signal pp_5_4 : std_logic;
signal pp_6_4 : std_logic;
signal pp_7_4 : std_logic;
signal pp_8_4 : std_logic;
signal pp_9_4 : std_logic;
signal pp_10_4 : std_logic;
signal pp_11_4 : std_logic;
signal pp_12_4 : std_logic;
signal pp_13_4 : std_logic;
signal pp_14_4 : std_logic;
signal pp_15_4 : std_logic;
signal pp_0_5 : std_logic;
signal pp_1_5 : std_logic;
signal pp_2_5 : std_logic;
signal pp_3_5 : std_logic;
signal pp_4_5 : std_logic;
signal pp_5_5 : std_logic;
signal pp_6_5 : std_logic;
signal pp_7_5 : std_logic;
signal pp_8_5 : std_logic;
signal pp_9_5 : std_logic;
signal pp_10_5 : std_logic;
signal pp_11_5 : std_logic;
signal pp_12_5 : std_logic;
signal pp_13_5 : std_logic;
signal pp_14_5 : std_logic;
signal pp_15_5 : std_logic;
signal pp_0_6 : std_logic;
signal pp_1_6 : std_logic;
signal pp_2_6 : std_logic;
signal pp_3_6 : std_logic;
signal pp_4_6 : std_logic;
signal pp_5_6 : std_logic;
signal pp_6_6 : std_logic;
signal pp_7_6 : std_logic;
signal pp_8_6 : std_logic;
signal pp_9_6 : std_logic;
signal pp_10_6 : std_logic;
signal pp_11_6 : std_logic;
signal pp_12_6 : std_logic;
signal pp_13_6 : std_logic;
signal pp_14_6 : std_logic;
signal pp_15_6 : std_logic;
signal pp_0_7 : std_logic;
signal pp_1_7 : std_logic;
signal pp_2_7 : std_logic;
signal pp_3_7 : std_logic;
signal pp_4_7 : std_logic;
signal pp_5_7 : std_logic;
signal pp_6_7 : std_logic;
signal pp_7_7 : std_logic;
signal pp_8_7 : std_logic;
signal pp_9_7 : std_logic;
signal pp_10_7 : std_logic;
signal pp_11_7 : std_logic;
signal pp_12_7 : std_logic;
signal pp_13_7 : std_logic;
signal pp_14_7 : std_logic;
signal pp_15_7 : std_logic;
signal pp_0_8 : std_logic;
signal pp_1_8 : std_logic;
signal pp_2_8 : std_logic;
signal pp_3_8 : std_logic;
signal pp_4_8 : std_logic;
signal pp_5_8 : std_logic;
signal pp_6_8 : std_logic;
signal pp_7_8 : std_logic;
signal pp_8_8 : std_logic;
signal pp_9_8 : std_logic;
signal pp_10_8 : std_logic;
signal pp_11_8 : std_logic;
signal pp_12_8 : std_logic;
signal pp_13_8 : std_logic;
signal pp_14_8 : std_logic;
signal pp_15_8 : std_logic;
signal pp_0_9 : std_logic;
signal pp_1_9 : std_logic;
signal pp_2_9 : std_logic;
signal pp_3_9 : std_logic;
signal pp_4_9 : std_logic;
signal pp_5_9 : std_logic;
signal pp_6_9 : std_logic;
signal pp_7_9 : std_logic;
signal pp_8_9 : std_logic;
signal pp_9_9 : std_logic;
signal pp_10_9 : std_logic;
signal pp_11_9 : std_logic;
signal pp_12_9 : std_logic;
signal pp_13_9 : std_logic;
signal pp_14_9 : std_logic;
signal pp_15_9 : std_logic;
signal pp_0_10 : std_logic;
signal pp_1_10 : std_logic;
signal pp_2_10 : std_logic;
signal pp_3_10 : std_logic;
signal pp_4_10 : std_logic;
signal pp_5_10 : std_logic;
signal pp_6_10 : std_logic;
signal pp_7_10 : std_logic;
signal pp_8_10 : std_logic;
signal pp_9_10 : std_logic;
signal pp_10_10 : std_logic;
signal pp_11_10 : std_logic;
signal pp_12_10 : std_logic;
signal pp_13_10 : std_logic;
signal pp_14_10 : std_logic;
signal pp_15_10 : std_logic;
signal pp_0_11 : std_logic;
signal pp_1_11 : std_logic;
signal pp_2_11 : std_logic;
signal pp_3_11 : std_logic;
signal pp_4_11 : std_logic;
signal pp_5_11 : std_logic;
signal pp_6_11 : std_logic;
signal pp_7_11 : std_logic;
signal pp_8_11 : std_logic;
signal pp_9_11 : std_logic;
signal pp_10_11 : std_logic;
signal pp_11_11 : std_logic;
signal pp_12_11 : std_logic;
signal pp_13_11 : std_logic;
signal pp_14_11 : std_logic;
signal pp_15_11 : std_logic;
signal pp_0_12 : std_logic;
signal pp_1_12 : std_logic;
signal pp_2_12 : std_logic;
signal pp_3_12 : std_logic;
signal pp_4_12 : std_logic;
signal pp_5_12 : std_logic;
signal pp_6_12 : std_logic;
signal pp_7_12 : std_logic;
signal pp_8_12 : std_logic;
signal pp_9_12 : std_logic;
signal pp_10_12 : std_logic;
signal pp_11_12 : std_logic;
signal pp_12_12 : std_logic;
signal pp_13_12 : std_logic;
signal pp_14_12 : std_logic;
signal pp_15_12 : std_logic;
signal pp_0_13 : std_logic;
signal pp_1_13 : std_logic;
signal pp_2_13 : std_logic;
signal pp_3_13 : std_logic;
signal pp_4_13 : std_logic;
signal pp_5_13 : std_logic;
signal pp_6_13 : std_logic;
signal pp_7_13 : std_logic;
signal pp_8_13 : std_logic;
signal pp_9_13 : std_logic;
signal pp_10_13 : std_logic;
signal pp_11_13 : std_logic;
signal pp_12_13 : std_logic;
signal pp_13_13 : std_logic;
signal pp_14_13 : std_logic;
signal pp_15_13 : std_logic;
signal pp_0_14 : std_logic;
signal pp_1_14 : std_logic;
signal pp_2_14 : std_logic;
signal pp_3_14 : std_logic;
signal pp_4_14 : std_logic;
signal pp_5_14 : std_logic;
signal pp_6_14 : std_logic;
signal pp_7_14 : std_logic;
signal pp_8_14 : std_logic;
signal pp_9_14 : std_logic;
signal pp_10_14 : std_logic;
signal pp_11_14 : std_logic;
signal pp_12_14 : std_logic;
signal pp_13_14 : std_logic;
signal pp_14_14 : std_logic;
signal pp_15_14 : std_logic;
signal pp_0_15 : std_logic;
signal pp_1_15 : std_logic;
signal pp_2_15 : std_logic;
signal pp_3_15 : std_logic;
signal pp_4_15 : std_logic;
signal pp_5_15 : std_logic;
signal pp_6_15 : std_logic;
signal pp_7_15 : std_logic;
signal pp_8_15 : std_logic;
signal pp_9_15 : std_logic;
signal pp_10_15 : std_logic;
signal pp_11_15 : std_logic;
signal pp_12_15 : std_logic;
signal pp_13_15 : std_logic;
signal pp_14_15 : std_logic;
signal pp_15_15 : std_logic;
signal ripple_carry_1 : std_logic;
signal ripple_carry_2 : std_logic;
signal ripple_carry_3 : std_logic;
signal ripple_carry_4 : std_logic;
signal ripple_carry_5 : std_logic;
signal ripple_carry_6 : std_logic;
signal ripple_carry_7 : std_logic;
signal ripple_carry_8 : std_logic;
signal ripple_carry_9 : std_logic;
signal ripple_carry_10 : std_logic;
signal ripple_carry_11 : std_logic;
signal ripple_carry_12 : std_logic;
signal ripple_carry_13 : std_logic;
signal ripple_carry_14 : std_logic;
signal ripple_carry_15 : std_logic;
signal ripple_carry_16 : std_logic;
signal ripple_carry_17 : std_logic;
signal ripple_carry_18 : std_logic;
signal ripple_carry_19 : std_logic;
signal ripple_carry_20 : std_logic;
signal ripple_carry_21 : std_logic;
signal ripple_carry_22 : std_logic;
signal ripple_carry_23 : std_logic;
signal ripple_carry_24 : std_logic;
signal ripple_carry_25 : std_logic;
signal ripple_carry_26 : std_logic;
signal ripple_carry_27 : std_logic;
signal ripple_carry_28 : std_logic;
signal ripple_carry_29 : std_logic;
signal ripple_carry_30 : std_logic;

begin

    
        half_adder_84639 : half_adder
            port map (
                a => pp_0_15,
                b => pp_1_14,
                s => sum_757675,
                Cout => cout_769389
            );
        

        half_adder_18278 : half_adder
            port map (
                a => pp_1_15,
                b => pp_2_14,
                s => sum_932346,
                Cout => cout_39739
            );
        

        full_adder_49951 : full_adder
            port map (
                a => sum_757675,
                b => pp_2_13,
                Cin => pp_3_12,
                s => sum_659249,
                Cout => cout_356642
            );
        

        full_adder_65933 : full_adder
            port map (
                a => sum_932346,
                b => cout_769389,
                Cin => pp_3_13,
                s => sum_47972,
                Cout => cout_39813
            );
        

        full_adder_50869 : full_adder
            port map (
                a => cout_39739,
                b => pp_2_15,
                Cin => pp_3_14,
                s => sum_753784,
                Cout => cout_172689
            );
        

        half_adder_38459 : half_adder
            port map (
                a => pp_0_14,
                b => pp_1_13,
                s => sum_754583,
                Cout => cout_624584
            );
        

        full_adder_29907 : full_adder
            port map (
                a => sum_754583,
                b => pp_2_12,
                Cin => pp_3_11,
                s => sum_538566,
                Cout => cout_172686
            );
        

        full_adder_34047 : full_adder
            port map (
                a => sum_659249,
                b => cout_624584,
                Cin => pp_4_11,
                s => sum_756610,
                Cout => cout_567486
            );
        

        full_adder_67817 : full_adder
            port map (
                a => sum_47972,
                b => cout_356642,
                Cin => pp_4_12,
                s => sum_914016,
                Cout => cout_913439
            );
        

        full_adder_44147 : full_adder
            port map (
                a => sum_753784,
                b => cout_39813,
                Cin => pp_4_13,
                s => sum_13181,
                Cout => cout_841917
            );
        

        full_adder_39753 : full_adder
            port map (
                a => cout_172689,
                b => pp_3_15,
                Cin => pp_4_14,
                s => sum_977726,
                Cout => cout_932234
            );
        

        half_adder_56721 : half_adder
            port map (
                a => pp_0_13,
                b => pp_1_12,
                s => sum_560320,
                Cout => cout_578344
            );
        

        full_adder_5591 : full_adder
            port map (
                a => sum_560320,
                b => pp_2_11,
                Cin => pp_3_10,
                s => sum_226390,
                Cout => cout_940010
            );
        

        full_adder_78010 : full_adder
            port map (
                a => sum_538566,
                b => cout_578344,
                Cin => pp_4_10,
                s => sum_766179,
                Cout => cout_491530
            );
        

        full_adder_77865 : full_adder
            port map (
                a => sum_756610,
                b => cout_172686,
                Cin => pp_5_10,
                s => sum_146247,
                Cout => cout_749783
            );
        

        full_adder_49099 : full_adder
            port map (
                a => sum_914016,
                b => cout_567486,
                Cin => pp_5_11,
                s => sum_722838,
                Cout => cout_905765
            );
        

        full_adder_76380 : full_adder
            port map (
                a => sum_13181,
                b => cout_913439,
                Cin => pp_5_12,
                s => sum_86012,
                Cout => cout_598245
            );
        

        full_adder_61456 : full_adder
            port map (
                a => sum_977726,
                b => cout_841917,
                Cin => pp_5_13,
                s => sum_492003,
                Cout => cout_191038
            );
        

        full_adder_3453 : full_adder
            port map (
                a => cout_932234,
                b => pp_4_15,
                Cin => pp_5_14,
                s => sum_618163,
                Cout => cout_578246
            );
        

        half_adder_25123 : half_adder
            port map (
                a => pp_0_12,
                b => pp_1_11,
                s => sum_910513,
                Cout => cout_94920
            );
        

        full_adder_1356 : full_adder
            port map (
                a => sum_910513,
                b => pp_2_10,
                Cin => pp_3_9,
                s => sum_990655,
                Cout => cout_976970
            );
        

        full_adder_59274 : full_adder
            port map (
                a => sum_226390,
                b => cout_94920,
                Cin => pp_4_9,
                s => sum_671502,
                Cout => cout_446076
            );
        

        full_adder_13211 : full_adder
            port map (
                a => sum_766179,
                b => cout_940010,
                Cin => pp_5_9,
                s => sum_411192,
                Cout => cout_461391
            );
        

        full_adder_32006 : full_adder
            port map (
                a => sum_146247,
                b => cout_491530,
                Cin => pp_6_9,
                s => sum_249416,
                Cout => cout_945951
            );
        

        full_adder_85363 : full_adder
            port map (
                a => sum_722838,
                b => cout_749783,
                Cin => pp_6_10,
                s => sum_686986,
                Cout => cout_712188
            );
        

        full_adder_64753 : full_adder
            port map (
                a => sum_86012,
                b => cout_905765,
                Cin => pp_6_11,
                s => sum_277628,
                Cout => cout_640546
            );
        

        full_adder_8933 : full_adder
            port map (
                a => sum_492003,
                b => cout_598245,
                Cin => pp_6_12,
                s => sum_287843,
                Cout => cout_275866
            );
        

        full_adder_72165 : full_adder
            port map (
                a => sum_618163,
                b => cout_191038,
                Cin => pp_6_13,
                s => sum_625716,
                Cout => cout_989486
            );
        

        full_adder_23342 : full_adder
            port map (
                a => cout_578246,
                b => pp_5_15,
                Cin => pp_6_14,
                s => sum_375464,
                Cout => cout_567696
            );
        

        half_adder_84703 : half_adder
            port map (
                a => pp_0_11,
                b => pp_1_10,
                s => sum_123741,
                Cout => cout_285703
            );
        

        full_adder_64591 : full_adder
            port map (
                a => sum_123741,
                b => pp_2_9,
                Cin => pp_3_8,
                s => sum_222046,
                Cout => cout_206738
            );
        

        full_adder_9428 : full_adder
            port map (
                a => sum_990655,
                b => cout_285703,
                Cin => pp_4_8,
                s => sum_7087,
                Cout => cout_262915
            );
        

        full_adder_74097 : full_adder
            port map (
                a => sum_671502,
                b => cout_976970,
                Cin => pp_5_8,
                s => sum_413141,
                Cout => cout_670764
            );
        

        full_adder_17995 : full_adder
            port map (
                a => sum_411192,
                b => cout_446076,
                Cin => pp_6_8,
                s => sum_380765,
                Cout => cout_918132
            );
        

        full_adder_40694 : full_adder
            port map (
                a => sum_249416,
                b => cout_461391,
                Cin => pp_7_8,
                s => sum_913153,
                Cout => cout_561087
            );
        

        full_adder_80896 : full_adder
            port map (
                a => sum_686986,
                b => cout_945951,
                Cin => pp_7_9,
                s => sum_390680,
                Cout => cout_357374
            );
        

        full_adder_69368 : full_adder
            port map (
                a => sum_277628,
                b => cout_712188,
                Cin => pp_7_10,
                s => sum_616616,
                Cout => cout_786530
            );
        

        full_adder_70736 : full_adder
            port map (
                a => sum_287843,
                b => cout_640546,
                Cin => pp_7_11,
                s => sum_863047,
                Cout => cout_960948
            );
        

        full_adder_32897 : full_adder
            port map (
                a => sum_625716,
                b => cout_275866,
                Cin => pp_7_12,
                s => sum_774946,
                Cout => cout_203266
            );
        

        full_adder_44913 : full_adder
            port map (
                a => sum_375464,
                b => cout_989486,
                Cin => pp_7_13,
                s => sum_961775,
                Cout => cout_860843
            );
        

        full_adder_71807 : full_adder
            port map (
                a => cout_567696,
                b => pp_6_15,
                Cin => pp_7_14,
                s => sum_451910,
                Cout => cout_420673
            );
        

        half_adder_92802 : half_adder
            port map (
                a => pp_0_10,
                b => pp_1_9,
                s => sum_327095,
                Cout => cout_863399
            );
        

        full_adder_54574 : full_adder
            port map (
                a => sum_327095,
                b => pp_2_8,
                Cin => pp_3_7,
                s => sum_274274,
                Cout => cout_930231
            );
        

        full_adder_22104 : full_adder
            port map (
                a => sum_222046,
                b => cout_863399,
                Cin => pp_4_7,
                s => sum_194968,
                Cout => cout_157897
            );
        

        full_adder_84059 : full_adder
            port map (
                a => sum_7087,
                b => cout_206738,
                Cin => pp_5_7,
                s => sum_24183,
                Cout => cout_551891
            );
        

        full_adder_67850 : full_adder
            port map (
                a => sum_413141,
                b => cout_262915,
                Cin => pp_6_7,
                s => sum_349866,
                Cout => cout_433248
            );
        

        full_adder_50768 : full_adder
            port map (
                a => sum_380765,
                b => cout_670764,
                Cin => pp_7_7,
                s => sum_797979,
                Cout => cout_187818
            );
        

        full_adder_61000 : full_adder
            port map (
                a => sum_913153,
                b => cout_918132,
                Cin => pp_8_7,
                s => sum_427572,
                Cout => cout_923055
            );
        

        full_adder_60253 : full_adder
            port map (
                a => sum_390680,
                b => cout_561087,
                Cin => pp_8_8,
                s => sum_797511,
                Cout => cout_878210
            );
        

        full_adder_14085 : full_adder
            port map (
                a => sum_616616,
                b => cout_357374,
                Cin => pp_8_9,
                s => sum_409507,
                Cout => cout_697098
            );
        

        full_adder_16784 : full_adder
            port map (
                a => sum_863047,
                b => cout_786530,
                Cin => pp_8_10,
                s => sum_181157,
                Cout => cout_537561
            );
        

        full_adder_20636 : full_adder
            port map (
                a => sum_774946,
                b => cout_960948,
                Cin => pp_8_11,
                s => sum_315286,
                Cout => cout_987740
            );
        

        full_adder_45141 : full_adder
            port map (
                a => sum_961775,
                b => cout_203266,
                Cin => pp_8_12,
                s => sum_404304,
                Cout => cout_22433
            );
        

        full_adder_4130 : full_adder
            port map (
                a => sum_451910,
                b => cout_860843,
                Cin => pp_8_13,
                s => sum_383733,
                Cout => cout_632990
            );
        

        full_adder_8096 : full_adder
            port map (
                a => cout_420673,
                b => pp_7_15,
                Cin => pp_8_14,
                s => sum_360115,
                Cout => cout_174525
            );
        

        half_adder_21996 : half_adder
            port map (
                a => pp_0_9,
                b => pp_1_8,
                s => sum_208632,
                Cout => cout_771281
            );
        

        full_adder_28476 : full_adder
            port map (
                a => sum_208632,
                b => pp_2_7,
                Cin => pp_3_6,
                s => sum_372567,
                Cout => cout_539978
            );
        

        full_adder_21468 : full_adder
            port map (
                a => sum_274274,
                b => cout_771281,
                Cin => pp_4_6,
                s => sum_246201,
                Cout => cout_258710
            );
        

        full_adder_66833 : full_adder
            port map (
                a => sum_194968,
                b => cout_930231,
                Cin => pp_5_6,
                s => sum_903520,
                Cout => cout_815001
            );
        

        full_adder_93690 : full_adder
            port map (
                a => sum_24183,
                b => cout_157897,
                Cin => pp_6_6,
                s => sum_774546,
                Cout => cout_346012
            );
        

        full_adder_34770 : full_adder
            port map (
                a => sum_349866,
                b => cout_551891,
                Cin => pp_7_6,
                s => sum_960667,
                Cout => cout_937613
            );
        

        full_adder_33603 : full_adder
            port map (
                a => sum_797979,
                b => cout_433248,
                Cin => pp_8_6,
                s => sum_705137,
                Cout => cout_153737
            );
        

        full_adder_91959 : full_adder
            port map (
                a => sum_427572,
                b => cout_187818,
                Cin => pp_9_6,
                s => sum_149238,
                Cout => cout_702253
            );
        

        full_adder_9885 : full_adder
            port map (
                a => sum_797511,
                b => cout_923055,
                Cin => pp_9_7,
                s => sum_388368,
                Cout => cout_529839
            );
        

        full_adder_12398 : full_adder
            port map (
                a => sum_409507,
                b => cout_878210,
                Cin => pp_9_8,
                s => sum_419352,
                Cout => cout_167953
            );
        

        full_adder_82673 : full_adder
            port map (
                a => sum_181157,
                b => cout_697098,
                Cin => pp_9_9,
                s => sum_796092,
                Cout => cout_759053
            );
        

        full_adder_47970 : full_adder
            port map (
                a => sum_315286,
                b => cout_537561,
                Cin => pp_9_10,
                s => sum_135226,
                Cout => cout_725574
            );
        

        full_adder_87409 : full_adder
            port map (
                a => sum_404304,
                b => cout_987740,
                Cin => pp_9_11,
                s => sum_165325,
                Cout => cout_242304
            );
        

        full_adder_93531 : full_adder
            port map (
                a => sum_383733,
                b => cout_22433,
                Cin => pp_9_12,
                s => sum_669906,
                Cout => cout_810450
            );
        

        full_adder_30513 : full_adder
            port map (
                a => sum_360115,
                b => cout_632990,
                Cin => pp_9_13,
                s => sum_711628,
                Cout => cout_666929
            );
        

        full_adder_87980 : full_adder
            port map (
                a => cout_174525,
                b => pp_8_15,
                Cin => pp_9_14,
                s => sum_410690,
                Cout => cout_22372
            );
        

        half_adder_57621 : half_adder
            port map (
                a => pp_0_8,
                b => pp_1_7,
                s => sum_230909,
                Cout => cout_727671
            );
        

        full_adder_68947 : full_adder
            port map (
                a => sum_230909,
                b => pp_2_6,
                Cin => pp_3_5,
                s => sum_905500,
                Cout => cout_525986
            );
        

        full_adder_7857 : full_adder
            port map (
                a => sum_372567,
                b => cout_727671,
                Cin => pp_4_5,
                s => sum_975960,
                Cout => cout_263090
            );
        

        full_adder_26221 : full_adder
            port map (
                a => sum_246201,
                b => cout_539978,
                Cin => pp_5_5,
                s => sum_21048,
                Cout => cout_649712
            );
        

        full_adder_16777 : full_adder
            port map (
                a => sum_903520,
                b => cout_258710,
                Cin => pp_6_5,
                s => sum_592564,
                Cout => cout_366028
            );
        

        full_adder_75262 : full_adder
            port map (
                a => sum_774546,
                b => cout_815001,
                Cin => pp_7_5,
                s => sum_272977,
                Cout => cout_69885
            );
        

        full_adder_41347 : full_adder
            port map (
                a => sum_960667,
                b => cout_346012,
                Cin => pp_8_5,
                s => sum_387065,
                Cout => cout_272868
            );
        

        full_adder_90273 : full_adder
            port map (
                a => sum_705137,
                b => cout_937613,
                Cin => pp_9_5,
                s => sum_182442,
                Cout => cout_922087
            );
        

        full_adder_74877 : full_adder
            port map (
                a => sum_149238,
                b => cout_153737,
                Cin => pp_10_5,
                s => sum_409,
                Cout => cout_821655
            );
        

        full_adder_41452 : full_adder
            port map (
                a => sum_388368,
                b => cout_702253,
                Cin => pp_10_6,
                s => sum_808671,
                Cout => cout_61302
            );
        

        full_adder_75412 : full_adder
            port map (
                a => sum_419352,
                b => cout_529839,
                Cin => pp_10_7,
                s => sum_113860,
                Cout => cout_327241
            );
        

        full_adder_27121 : full_adder
            port map (
                a => sum_796092,
                b => cout_167953,
                Cin => pp_10_8,
                s => sum_248889,
                Cout => cout_82325
            );
        

        full_adder_53236 : full_adder
            port map (
                a => sum_135226,
                b => cout_759053,
                Cin => pp_10_9,
                s => sum_343072,
                Cout => cout_791728
            );
        

        full_adder_37334 : full_adder
            port map (
                a => sum_165325,
                b => cout_725574,
                Cin => pp_10_10,
                s => sum_659836,
                Cout => cout_684959
            );
        

        full_adder_76637 : full_adder
            port map (
                a => sum_669906,
                b => cout_242304,
                Cin => pp_10_11,
                s => sum_658736,
                Cout => cout_846804
            );
        

        full_adder_16642 : full_adder
            port map (
                a => sum_711628,
                b => cout_810450,
                Cin => pp_10_12,
                s => sum_241703,
                Cout => cout_974942
            );
        

        full_adder_7188 : full_adder
            port map (
                a => sum_410690,
                b => cout_666929,
                Cin => pp_10_13,
                s => sum_324032,
                Cout => cout_889121
            );
        

        full_adder_65228 : full_adder
            port map (
                a => cout_22372,
                b => pp_9_15,
                Cin => pp_10_14,
                s => sum_647575,
                Cout => cout_904012
            );
        

        half_adder_1679 : half_adder
            port map (
                a => pp_0_7,
                b => pp_1_6,
                s => sum_310349,
                Cout => cout_82769
            );
        

        full_adder_66587 : full_adder
            port map (
                a => sum_310349,
                b => pp_2_5,
                Cin => pp_3_4,
                s => sum_641583,
                Cout => cout_199542
            );
        

        full_adder_63541 : full_adder
            port map (
                a => sum_905500,
                b => cout_82769,
                Cin => pp_4_4,
                s => sum_752893,
                Cout => cout_936261
            );
        

        full_adder_87000 : full_adder
            port map (
                a => sum_975960,
                b => cout_525986,
                Cin => pp_5_4,
                s => sum_548921,
                Cout => cout_138274
            );
        

        full_adder_15465 : full_adder
            port map (
                a => sum_21048,
                b => cout_263090,
                Cin => pp_6_4,
                s => sum_461182,
                Cout => cout_599211
            );
        

        full_adder_62439 : full_adder
            port map (
                a => sum_592564,
                b => cout_649712,
                Cin => pp_7_4,
                s => sum_319630,
                Cout => cout_152176
            );
        

        full_adder_24145 : full_adder
            port map (
                a => sum_272977,
                b => cout_366028,
                Cin => pp_8_4,
                s => sum_533069,
                Cout => cout_111262
            );
        

        full_adder_44450 : full_adder
            port map (
                a => sum_387065,
                b => cout_69885,
                Cin => pp_9_4,
                s => sum_887964,
                Cout => cout_284285
            );
        

        full_adder_14038 : full_adder
            port map (
                a => sum_182442,
                b => cout_272868,
                Cin => pp_10_4,
                s => sum_835449,
                Cout => cout_139640
            );
        

        full_adder_63826 : full_adder
            port map (
                a => sum_409,
                b => cout_922087,
                Cin => pp_11_4,
                s => sum_993754,
                Cout => cout_177382
            );
        

        full_adder_92373 : full_adder
            port map (
                a => sum_808671,
                b => cout_821655,
                Cin => pp_11_5,
                s => sum_504281,
                Cout => cout_5038
            );
        

        full_adder_84399 : full_adder
            port map (
                a => sum_113860,
                b => cout_61302,
                Cin => pp_11_6,
                s => sum_909922,
                Cout => cout_662043
            );
        

        full_adder_83256 : full_adder
            port map (
                a => sum_248889,
                b => cout_327241,
                Cin => pp_11_7,
                s => sum_766402,
                Cout => cout_63167
            );
        

        full_adder_44438 : full_adder
            port map (
                a => sum_343072,
                b => cout_82325,
                Cin => pp_11_8,
                s => sum_439931,
                Cout => cout_599694
            );
        

        full_adder_20123 : full_adder
            port map (
                a => sum_659836,
                b => cout_791728,
                Cin => pp_11_9,
                s => sum_911256,
                Cout => cout_952902
            );
        

        full_adder_27557 : full_adder
            port map (
                a => sum_658736,
                b => cout_684959,
                Cin => pp_11_10,
                s => sum_530689,
                Cout => cout_606994
            );
        

        full_adder_9258 : full_adder
            port map (
                a => sum_241703,
                b => cout_846804,
                Cin => pp_11_11,
                s => sum_442354,
                Cout => cout_738496
            );
        

        full_adder_12555 : full_adder
            port map (
                a => sum_324032,
                b => cout_974942,
                Cin => pp_11_12,
                s => sum_85078,
                Cout => cout_43875
            );
        

        full_adder_31125 : full_adder
            port map (
                a => sum_647575,
                b => cout_889121,
                Cin => pp_11_13,
                s => sum_716697,
                Cout => cout_180198
            );
        

        full_adder_95749 : full_adder
            port map (
                a => cout_904012,
                b => pp_10_15,
                Cin => pp_11_14,
                s => sum_579393,
                Cout => cout_401825
            );
        

        half_adder_16747 : half_adder
            port map (
                a => pp_0_6,
                b => pp_1_5,
                s => sum_742414,
                Cout => cout_276204
            );
        

        full_adder_39175 : full_adder
            port map (
                a => sum_742414,
                b => pp_2_4,
                Cin => pp_3_3,
                s => sum_878840,
                Cout => cout_413325
            );
        

        full_adder_56293 : full_adder
            port map (
                a => sum_641583,
                b => cout_276204,
                Cin => pp_4_3,
                s => sum_952338,
                Cout => cout_227086
            );
        

        full_adder_61251 : full_adder
            port map (
                a => sum_752893,
                b => cout_199542,
                Cin => pp_5_3,
                s => sum_922115,
                Cout => cout_232219
            );
        

        full_adder_58713 : full_adder
            port map (
                a => sum_548921,
                b => cout_936261,
                Cin => pp_6_3,
                s => sum_584013,
                Cout => cout_403061
            );
        

        full_adder_6407 : full_adder
            port map (
                a => sum_461182,
                b => cout_138274,
                Cin => pp_7_3,
                s => sum_859480,
                Cout => cout_928577
            );
        

        full_adder_1025 : full_adder
            port map (
                a => sum_319630,
                b => cout_599211,
                Cin => pp_8_3,
                s => sum_807794,
                Cout => cout_847359
            );
        

        full_adder_15609 : full_adder
            port map (
                a => sum_533069,
                b => cout_152176,
                Cin => pp_9_3,
                s => sum_202927,
                Cout => cout_299193
            );
        

        full_adder_24147 : full_adder
            port map (
                a => sum_887964,
                b => cout_111262,
                Cin => pp_10_3,
                s => sum_830004,
                Cout => cout_599178
            );
        

        full_adder_90828 : full_adder
            port map (
                a => sum_835449,
                b => cout_284285,
                Cin => pp_11_3,
                s => sum_418595,
                Cout => cout_717070
            );
        

        full_adder_18538 : full_adder
            port map (
                a => sum_993754,
                b => cout_139640,
                Cin => pp_12_3,
                s => sum_877555,
                Cout => cout_186640
            );
        

        full_adder_77591 : full_adder
            port map (
                a => sum_504281,
                b => cout_177382,
                Cin => pp_12_4,
                s => sum_885640,
                Cout => cout_744469
            );
        

        full_adder_30082 : full_adder
            port map (
                a => sum_909922,
                b => cout_5038,
                Cin => pp_12_5,
                s => sum_568950,
                Cout => cout_217500
            );
        

        full_adder_38481 : full_adder
            port map (
                a => sum_766402,
                b => cout_662043,
                Cin => pp_12_6,
                s => sum_37576,
                Cout => cout_543060
            );
        

        full_adder_20555 : full_adder
            port map (
                a => sum_439931,
                b => cout_63167,
                Cin => pp_12_7,
                s => sum_871425,
                Cout => cout_380034
            );
        

        full_adder_4479 : full_adder
            port map (
                a => sum_911256,
                b => cout_599694,
                Cin => pp_12_8,
                s => sum_963006,
                Cout => cout_960555
            );
        

        full_adder_64588 : full_adder
            port map (
                a => sum_530689,
                b => cout_952902,
                Cin => pp_12_9,
                s => sum_179806,
                Cout => cout_909674
            );
        

        full_adder_60286 : full_adder
            port map (
                a => sum_442354,
                b => cout_606994,
                Cin => pp_12_10,
                s => sum_622556,
                Cout => cout_6366
            );
        

        full_adder_53515 : full_adder
            port map (
                a => sum_85078,
                b => cout_738496,
                Cin => pp_12_11,
                s => sum_100853,
                Cout => cout_241998
            );
        

        full_adder_65697 : full_adder
            port map (
                a => sum_716697,
                b => cout_43875,
                Cin => pp_12_12,
                s => sum_590812,
                Cout => cout_189105
            );
        

        full_adder_16870 : full_adder
            port map (
                a => sum_579393,
                b => cout_180198,
                Cin => pp_12_13,
                s => sum_853972,
                Cout => cout_908865
            );
        

        full_adder_60841 : full_adder
            port map (
                a => cout_401825,
                b => pp_11_15,
                Cin => pp_12_14,
                s => sum_487151,
                Cout => cout_428500
            );
        

        half_adder_64930 : half_adder
            port map (
                a => pp_0_5,
                b => pp_1_4,
                s => sum_964352,
                Cout => cout_5705
            );
        

        full_adder_49224 : full_adder
            port map (
                a => sum_964352,
                b => pp_2_3,
                Cin => pp_3_2,
                s => sum_190083,
                Cout => cout_44270
            );
        

        full_adder_66590 : full_adder
            port map (
                a => sum_878840,
                b => cout_5705,
                Cin => pp_4_2,
                s => sum_155461,
                Cout => cout_752478
            );
        

        full_adder_15706 : full_adder
            port map (
                a => sum_952338,
                b => cout_413325,
                Cin => pp_5_2,
                s => sum_70271,
                Cout => cout_103199
            );
        

        full_adder_59520 : full_adder
            port map (
                a => sum_922115,
                b => cout_227086,
                Cin => pp_6_2,
                s => sum_325561,
                Cout => cout_503461
            );
        

        full_adder_74757 : full_adder
            port map (
                a => sum_584013,
                b => cout_232219,
                Cin => pp_7_2,
                s => sum_384618,
                Cout => cout_554463
            );
        

        full_adder_77238 : full_adder
            port map (
                a => sum_859480,
                b => cout_403061,
                Cin => pp_8_2,
                s => sum_610884,
                Cout => cout_963328
            );
        

        full_adder_72679 : full_adder
            port map (
                a => sum_807794,
                b => cout_928577,
                Cin => pp_9_2,
                s => sum_527017,
                Cout => cout_836750
            );
        

        full_adder_9505 : full_adder
            port map (
                a => sum_202927,
                b => cout_847359,
                Cin => pp_10_2,
                s => sum_330037,
                Cout => cout_845115
            );
        

        full_adder_94072 : full_adder
            port map (
                a => sum_830004,
                b => cout_299193,
                Cin => pp_11_2,
                s => sum_617507,
                Cout => cout_187919
            );
        

        full_adder_4868 : full_adder
            port map (
                a => sum_418595,
                b => cout_599178,
                Cin => pp_12_2,
                s => sum_745173,
                Cout => cout_903116
            );
        

        full_adder_31188 : full_adder
            port map (
                a => sum_877555,
                b => cout_717070,
                Cin => pp_13_2,
                s => sum_107552,
                Cout => cout_57875
            );
        

        full_adder_68660 : full_adder
            port map (
                a => sum_885640,
                b => cout_186640,
                Cin => pp_13_3,
                s => sum_3669,
                Cout => cout_924814
            );
        

        full_adder_79547 : full_adder
            port map (
                a => sum_568950,
                b => cout_744469,
                Cin => pp_13_4,
                s => sum_890133,
                Cout => cout_752540
            );
        

        full_adder_16834 : full_adder
            port map (
                a => sum_37576,
                b => cout_217500,
                Cin => pp_13_5,
                s => sum_285660,
                Cout => cout_750878
            );
        

        full_adder_47670 : full_adder
            port map (
                a => sum_871425,
                b => cout_543060,
                Cin => pp_13_6,
                s => sum_865435,
                Cout => cout_347189
            );
        

        full_adder_47871 : full_adder
            port map (
                a => sum_963006,
                b => cout_380034,
                Cin => pp_13_7,
                s => sum_165169,
                Cout => cout_903701
            );
        

        full_adder_68974 : full_adder
            port map (
                a => sum_179806,
                b => cout_960555,
                Cin => pp_13_8,
                s => sum_161296,
                Cout => cout_9966
            );
        

        full_adder_68218 : full_adder
            port map (
                a => sum_622556,
                b => cout_909674,
                Cin => pp_13_9,
                s => sum_210485,
                Cout => cout_154367
            );
        

        full_adder_82864 : full_adder
            port map (
                a => sum_100853,
                b => cout_6366,
                Cin => pp_13_10,
                s => sum_940061,
                Cout => cout_777808
            );
        

        full_adder_16360 : full_adder
            port map (
                a => sum_590812,
                b => cout_241998,
                Cin => pp_13_11,
                s => sum_556282,
                Cout => cout_918370
            );
        

        full_adder_90077 : full_adder
            port map (
                a => sum_853972,
                b => cout_189105,
                Cin => pp_13_12,
                s => sum_409267,
                Cout => cout_765436
            );
        

        full_adder_53568 : full_adder
            port map (
                a => sum_487151,
                b => cout_908865,
                Cin => pp_13_13,
                s => sum_16716,
                Cout => cout_743533
            );
        

        full_adder_94586 : full_adder
            port map (
                a => cout_428500,
                b => pp_12_15,
                Cin => pp_13_14,
                s => sum_128628,
                Cout => cout_809894
            );
        

        half_adder_63696 : half_adder
            port map (
                a => pp_0_4,
                b => pp_1_3,
                s => sum_151833,
                Cout => cout_442253
            );
        

        full_adder_52824 : full_adder
            port map (
                a => sum_151833,
                b => pp_2_2,
                Cin => pp_3_1,
                s => sum_491221,
                Cout => cout_681963
            );
        

        full_adder_22162 : full_adder
            port map (
                a => sum_190083,
                b => cout_442253,
                Cin => pp_4_1,
                s => sum_372577,
                Cout => cout_12222
            );
        

        full_adder_49603 : full_adder
            port map (
                a => sum_155461,
                b => cout_44270,
                Cin => pp_5_1,
                s => sum_352335,
                Cout => cout_194219
            );
        

        full_adder_24789 : full_adder
            port map (
                a => sum_70271,
                b => cout_752478,
                Cin => pp_6_1,
                s => sum_218632,
                Cout => cout_283181
            );
        

        full_adder_93689 : full_adder
            port map (
                a => sum_325561,
                b => cout_103199,
                Cin => pp_7_1,
                s => sum_509457,
                Cout => cout_801902
            );
        

        full_adder_72712 : full_adder
            port map (
                a => sum_384618,
                b => cout_503461,
                Cin => pp_8_1,
                s => sum_813250,
                Cout => cout_597879
            );
        

        full_adder_87804 : full_adder
            port map (
                a => sum_610884,
                b => cout_554463,
                Cin => pp_9_1,
                s => sum_436895,
                Cout => cout_52308
            );
        

        full_adder_58753 : full_adder
            port map (
                a => sum_527017,
                b => cout_963328,
                Cin => pp_10_1,
                s => sum_608641,
                Cout => cout_230642
            );
        

        full_adder_69463 : full_adder
            port map (
                a => sum_330037,
                b => cout_836750,
                Cin => pp_11_1,
                s => sum_75594,
                Cout => cout_269720
            );
        

        full_adder_7886 : full_adder
            port map (
                a => sum_617507,
                b => cout_845115,
                Cin => pp_12_1,
                s => sum_538112,
                Cout => cout_612378
            );
        

        full_adder_7163 : full_adder
            port map (
                a => sum_745173,
                b => cout_187919,
                Cin => pp_13_1,
                s => sum_752554,
                Cout => cout_390278
            );
        

        full_adder_62881 : full_adder
            port map (
                a => sum_107552,
                b => cout_903116,
                Cin => pp_14_1,
                s => sum_447835,
                Cout => cout_81863
            );
        

        full_adder_12381 : full_adder
            port map (
                a => sum_3669,
                b => cout_57875,
                Cin => pp_14_2,
                s => sum_604064,
                Cout => cout_665374
            );
        

        full_adder_75297 : full_adder
            port map (
                a => sum_890133,
                b => cout_924814,
                Cin => pp_14_3,
                s => sum_602802,
                Cout => cout_313284
            );
        

        full_adder_77296 : full_adder
            port map (
                a => sum_285660,
                b => cout_752540,
                Cin => pp_14_4,
                s => sum_447776,
                Cout => cout_610447
            );
        

        full_adder_56975 : full_adder
            port map (
                a => sum_865435,
                b => cout_750878,
                Cin => pp_14_5,
                s => sum_846479,
                Cout => cout_58374
            );
        

        full_adder_81955 : full_adder
            port map (
                a => sum_165169,
                b => cout_347189,
                Cin => pp_14_6,
                s => sum_175238,
                Cout => cout_352004
            );
        

        full_adder_48637 : full_adder
            port map (
                a => sum_161296,
                b => cout_903701,
                Cin => pp_14_7,
                s => sum_101042,
                Cout => cout_120477
            );
        

        full_adder_5618 : full_adder
            port map (
                a => sum_210485,
                b => cout_9966,
                Cin => pp_14_8,
                s => sum_863612,
                Cout => cout_621744
            );
        

        full_adder_52142 : full_adder
            port map (
                a => sum_940061,
                b => cout_154367,
                Cin => pp_14_9,
                s => sum_292728,
                Cout => cout_253376
            );
        

        full_adder_9487 : full_adder
            port map (
                a => sum_556282,
                b => cout_777808,
                Cin => pp_14_10,
                s => sum_36423,
                Cout => cout_986139
            );
        

        full_adder_6558 : full_adder
            port map (
                a => sum_409267,
                b => cout_918370,
                Cin => pp_14_11,
                s => sum_763057,
                Cout => cout_830405
            );
        

        full_adder_84351 : full_adder
            port map (
                a => sum_16716,
                b => cout_765436,
                Cin => pp_14_12,
                s => sum_677725,
                Cout => cout_225273
            );
        

        full_adder_47334 : full_adder
            port map (
                a => sum_128628,
                b => cout_743533,
                Cin => pp_14_13,
                s => sum_924856,
                Cout => cout_105480
            );
        

        full_adder_59158 : full_adder
            port map (
                a => cout_809894,
                b => pp_13_15,
                Cin => pp_14_14,
                s => sum_653807,
                Cout => cout_683444
            );
        

        half_adder_73637 : half_adder
            port map (
                a => pp_0_3,
                b => pp_1_2,
                s => sum_393354,
                Cout => cout_773384
            );
        

        full_adder_42305 : full_adder
            port map (
                a => sum_393354,
                b => pp_2_1,
                Cin => pp_3_0,
                s => sum_454017,
                Cout => cout_648852
            );
        

        full_adder_9911 : full_adder
            port map (
                a => sum_491221,
                b => cout_773384,
                Cin => pp_4_0,
                s => sum_615388,
                Cout => cout_622190
            );
        

        full_adder_60996 : full_adder
            port map (
                a => sum_372577,
                b => cout_681963,
                Cin => pp_5_0,
                s => sum_307052,
                Cout => cout_296984
            );
        

        full_adder_56682 : full_adder
            port map (
                a => sum_352335,
                b => cout_12222,
                Cin => pp_6_0,
                s => sum_957721,
                Cout => cout_372708
            );
        

        full_adder_852 : full_adder
            port map (
                a => sum_218632,
                b => cout_194219,
                Cin => pp_7_0,
                s => sum_910907,
                Cout => cout_87182
            );
        

        full_adder_53946 : full_adder
            port map (
                a => sum_509457,
                b => cout_283181,
                Cin => pp_8_0,
                s => sum_190554,
                Cout => cout_901791
            );
        

        full_adder_94055 : full_adder
            port map (
                a => sum_813250,
                b => cout_801902,
                Cin => pp_9_0,
                s => sum_108552,
                Cout => cout_938354
            );
        

        full_adder_13911 : full_adder
            port map (
                a => sum_436895,
                b => cout_597879,
                Cin => pp_10_0,
                s => sum_871398,
                Cout => cout_899840
            );
        

        full_adder_81279 : full_adder
            port map (
                a => sum_608641,
                b => cout_52308,
                Cin => pp_11_0,
                s => sum_748543,
                Cout => cout_473235
            );
        

        full_adder_81843 : full_adder
            port map (
                a => sum_75594,
                b => cout_230642,
                Cin => pp_12_0,
                s => sum_620884,
                Cout => cout_502572
            );
        

        full_adder_64886 : full_adder
            port map (
                a => sum_538112,
                b => cout_269720,
                Cin => pp_13_0,
                s => sum_835826,
                Cout => cout_615799
            );
        

        full_adder_84248 : full_adder
            port map (
                a => sum_752554,
                b => cout_612378,
                Cin => pp_14_0,
                s => sum_747437,
                Cout => cout_907232
            );
        

        full_adder_18298 : full_adder
            port map (
                a => sum_447835,
                b => cout_390278,
                Cin => pp_15_0,
                s => sum_408519,
                Cout => cout_273843
            );
        

        full_adder_69625 : full_adder
            port map (
                a => sum_604064,
                b => cout_81863,
                Cin => pp_15_1,
                s => sum_825709,
                Cout => cout_593623
            );
        

        full_adder_94627 : full_adder
            port map (
                a => sum_602802,
                b => cout_665374,
                Cin => pp_15_2,
                s => sum_751602,
                Cout => cout_860894
            );
        

        full_adder_4131 : full_adder
            port map (
                a => sum_447776,
                b => cout_313284,
                Cin => pp_15_3,
                s => sum_739794,
                Cout => cout_336777
            );
        

        full_adder_52097 : full_adder
            port map (
                a => sum_846479,
                b => cout_610447,
                Cin => pp_15_4,
                s => sum_422751,
                Cout => cout_174675
            );
        

        full_adder_6319 : full_adder
            port map (
                a => sum_175238,
                b => cout_58374,
                Cin => pp_15_5,
                s => sum_573526,
                Cout => cout_622573
            );
        

        full_adder_28628 : full_adder
            port map (
                a => sum_101042,
                b => cout_352004,
                Cin => pp_15_6,
                s => sum_334672,
                Cout => cout_614796
            );
        

        full_adder_6375 : full_adder
            port map (
                a => sum_863612,
                b => cout_120477,
                Cin => pp_15_7,
                s => sum_445479,
                Cout => cout_694665
            );
        

        full_adder_56916 : full_adder
            port map (
                a => sum_292728,
                b => cout_621744,
                Cin => pp_15_8,
                s => sum_873056,
                Cout => cout_34362
            );
        

        full_adder_24330 : full_adder
            port map (
                a => sum_36423,
                b => cout_253376,
                Cin => pp_15_9,
                s => sum_860833,
                Cout => cout_288058
            );
        

        full_adder_38623 : full_adder
            port map (
                a => sum_763057,
                b => cout_986139,
                Cin => pp_15_10,
                s => sum_906512,
                Cout => cout_430498
            );
        

        full_adder_11222 : full_adder
            port map (
                a => sum_677725,
                b => cout_830405,
                Cin => pp_15_11,
                s => sum_319921,
                Cout => cout_310125
            );
        

        full_adder_76348 : full_adder
            port map (
                a => sum_924856,
                b => cout_225273,
                Cin => pp_15_12,
                s => sum_777791,
                Cout => cout_278529
            );
        

        full_adder_71974 : full_adder
            port map (
                a => sum_653807,
                b => cout_105480,
                Cin => pp_15_13,
                s => sum_134521,
                Cout => cout_907380
            );
        

        full_adder_89134 : full_adder
            port map (
                a => cout_683444,
                b => pp_14_15,
                Cin => pp_15_14,
                s => sum_453295,
                Cout => cout_505573
            );
        

        half_adder_96767 : half_adder
            port map (
                a => pp_0_2,
                b => pp_1_1,
                s => sum_652062,
                Cout => cout_734723
            );
        

        pp_0_0 <= a(0) and b(0);
        

        pp_1_0 <= a(1) and b(0);
        

        pp_2_0 <= a(2) and b(0);
        

        pp_3_0 <= a(3) and b(0);
        

        pp_4_0 <= a(4) and b(0);
        

        pp_5_0 <= a(5) and b(0);
        

        pp_6_0 <= a(6) and b(0);
        

        pp_7_0 <= a(7) and b(0);
        

        pp_8_0 <= a(8) and b(0);
        

        pp_9_0 <= a(9) and b(0);
        

        pp_10_0 <= a(10) and b(0);
        

        pp_11_0 <= a(11) and b(0);
        

        pp_12_0 <= a(12) and b(0);
        

        pp_13_0 <= a(13) and b(0);
        

        pp_14_0 <= a(14) and b(0);
        

        pp_15_0 <= a(15) and b(0);
        

        pp_0_1 <= a(0) and b(1);
        

        pp_1_1 <= a(1) and b(1);
        

        pp_2_1 <= a(2) and b(1);
        

        pp_3_1 <= a(3) and b(1);
        

        pp_4_1 <= a(4) and b(1);
        

        pp_5_1 <= a(5) and b(1);
        

        pp_6_1 <= a(6) and b(1);
        

        pp_7_1 <= a(7) and b(1);
        

        pp_8_1 <= a(8) and b(1);
        

        pp_9_1 <= a(9) and b(1);
        

        pp_10_1 <= a(10) and b(1);
        

        pp_11_1 <= a(11) and b(1);
        

        pp_12_1 <= a(12) and b(1);
        

        pp_13_1 <= a(13) and b(1);
        

        pp_14_1 <= a(14) and b(1);
        

        pp_15_1 <= a(15) and b(1);
        

        pp_0_2 <= a(0) and b(2);
        

        pp_1_2 <= a(1) and b(2);
        

        pp_2_2 <= a(2) and b(2);
        

        pp_3_2 <= a(3) and b(2);
        

        pp_4_2 <= a(4) and b(2);
        

        pp_5_2 <= a(5) and b(2);
        

        pp_6_2 <= a(6) and b(2);
        

        pp_7_2 <= a(7) and b(2);
        

        pp_8_2 <= a(8) and b(2);
        

        pp_9_2 <= a(9) and b(2);
        

        pp_10_2 <= a(10) and b(2);
        

        pp_11_2 <= a(11) and b(2);
        

        pp_12_2 <= a(12) and b(2);
        

        pp_13_2 <= a(13) and b(2);
        

        pp_14_2 <= a(14) and b(2);
        

        pp_15_2 <= a(15) and b(2);
        

        pp_0_3 <= a(0) and b(3);
        

        pp_1_3 <= a(1) and b(3);
        

        pp_2_3 <= a(2) and b(3);
        

        pp_3_3 <= a(3) and b(3);
        

        pp_4_3 <= a(4) and b(3);
        

        pp_5_3 <= a(5) and b(3);
        

        pp_6_3 <= a(6) and b(3);
        

        pp_7_3 <= a(7) and b(3);
        

        pp_8_3 <= a(8) and b(3);
        

        pp_9_3 <= a(9) and b(3);
        

        pp_10_3 <= a(10) and b(3);
        

        pp_11_3 <= a(11) and b(3);
        

        pp_12_3 <= a(12) and b(3);
        

        pp_13_3 <= a(13) and b(3);
        

        pp_14_3 <= a(14) and b(3);
        

        pp_15_3 <= a(15) and b(3);
        

        pp_0_4 <= a(0) and b(4);
        

        pp_1_4 <= a(1) and b(4);
        

        pp_2_4 <= a(2) and b(4);
        

        pp_3_4 <= a(3) and b(4);
        

        pp_4_4 <= a(4) and b(4);
        

        pp_5_4 <= a(5) and b(4);
        

        pp_6_4 <= a(6) and b(4);
        

        pp_7_4 <= a(7) and b(4);
        

        pp_8_4 <= a(8) and b(4);
        

        pp_9_4 <= a(9) and b(4);
        

        pp_10_4 <= a(10) and b(4);
        

        pp_11_4 <= a(11) and b(4);
        

        pp_12_4 <= a(12) and b(4);
        

        pp_13_4 <= a(13) and b(4);
        

        pp_14_4 <= a(14) and b(4);
        

        pp_15_4 <= a(15) and b(4);
        

        pp_0_5 <= a(0) and b(5);
        

        pp_1_5 <= a(1) and b(5);
        

        pp_2_5 <= a(2) and b(5);
        

        pp_3_5 <= a(3) and b(5);
        

        pp_4_5 <= a(4) and b(5);
        

        pp_5_5 <= a(5) and b(5);
        

        pp_6_5 <= a(6) and b(5);
        

        pp_7_5 <= a(7) and b(5);
        

        pp_8_5 <= a(8) and b(5);
        

        pp_9_5 <= a(9) and b(5);
        

        pp_10_5 <= a(10) and b(5);
        

        pp_11_5 <= a(11) and b(5);
        

        pp_12_5 <= a(12) and b(5);
        

        pp_13_5 <= a(13) and b(5);
        

        pp_14_5 <= a(14) and b(5);
        

        pp_15_5 <= a(15) and b(5);
        

        pp_0_6 <= a(0) and b(6);
        

        pp_1_6 <= a(1) and b(6);
        

        pp_2_6 <= a(2) and b(6);
        

        pp_3_6 <= a(3) and b(6);
        

        pp_4_6 <= a(4) and b(6);
        

        pp_5_6 <= a(5) and b(6);
        

        pp_6_6 <= a(6) and b(6);
        

        pp_7_6 <= a(7) and b(6);
        

        pp_8_6 <= a(8) and b(6);
        

        pp_9_6 <= a(9) and b(6);
        

        pp_10_6 <= a(10) and b(6);
        

        pp_11_6 <= a(11) and b(6);
        

        pp_12_6 <= a(12) and b(6);
        

        pp_13_6 <= a(13) and b(6);
        

        pp_14_6 <= a(14) and b(6);
        

        pp_15_6 <= a(15) and b(6);
        

        pp_0_7 <= a(0) and b(7);
        

        pp_1_7 <= a(1) and b(7);
        

        pp_2_7 <= a(2) and b(7);
        

        pp_3_7 <= a(3) and b(7);
        

        pp_4_7 <= a(4) and b(7);
        

        pp_5_7 <= a(5) and b(7);
        

        pp_6_7 <= a(6) and b(7);
        

        pp_7_7 <= a(7) and b(7);
        

        pp_8_7 <= a(8) and b(7);
        

        pp_9_7 <= a(9) and b(7);
        

        pp_10_7 <= a(10) and b(7);
        

        pp_11_7 <= a(11) and b(7);
        

        pp_12_7 <= a(12) and b(7);
        

        pp_13_7 <= a(13) and b(7);
        

        pp_14_7 <= a(14) and b(7);
        

        pp_15_7 <= a(15) and b(7);
        

        pp_0_8 <= a(0) and b(8);
        

        pp_1_8 <= a(1) and b(8);
        

        pp_2_8 <= a(2) and b(8);
        

        pp_3_8 <= a(3) and b(8);
        

        pp_4_8 <= a(4) and b(8);
        

        pp_5_8 <= a(5) and b(8);
        

        pp_6_8 <= a(6) and b(8);
        

        pp_7_8 <= a(7) and b(8);
        

        pp_8_8 <= a(8) and b(8);
        

        pp_9_8 <= a(9) and b(8);
        

        pp_10_8 <= a(10) and b(8);
        

        pp_11_8 <= a(11) and b(8);
        

        pp_12_8 <= a(12) and b(8);
        

        pp_13_8 <= a(13) and b(8);
        

        pp_14_8 <= a(14) and b(8);
        

        pp_15_8 <= a(15) and b(8);
        

        pp_0_9 <= a(0) and b(9);
        

        pp_1_9 <= a(1) and b(9);
        

        pp_2_9 <= a(2) and b(9);
        

        pp_3_9 <= a(3) and b(9);
        

        pp_4_9 <= a(4) and b(9);
        

        pp_5_9 <= a(5) and b(9);
        

        pp_6_9 <= a(6) and b(9);
        

        pp_7_9 <= a(7) and b(9);
        

        pp_8_9 <= a(8) and b(9);
        

        pp_9_9 <= a(9) and b(9);
        

        pp_10_9 <= a(10) and b(9);
        

        pp_11_9 <= a(11) and b(9);
        

        pp_12_9 <= a(12) and b(9);
        

        pp_13_9 <= a(13) and b(9);
        

        pp_14_9 <= a(14) and b(9);
        

        pp_15_9 <= a(15) and b(9);
        

        pp_0_10 <= a(0) and b(10);
        

        pp_1_10 <= a(1) and b(10);
        

        pp_2_10 <= a(2) and b(10);
        

        pp_3_10 <= a(3) and b(10);
        

        pp_4_10 <= a(4) and b(10);
        

        pp_5_10 <= a(5) and b(10);
        

        pp_6_10 <= a(6) and b(10);
        

        pp_7_10 <= a(7) and b(10);
        

        pp_8_10 <= a(8) and b(10);
        

        pp_9_10 <= a(9) and b(10);
        

        pp_10_10 <= a(10) and b(10);
        

        pp_11_10 <= a(11) and b(10);
        

        pp_12_10 <= a(12) and b(10);
        

        pp_13_10 <= a(13) and b(10);
        

        pp_14_10 <= a(14) and b(10);
        

        pp_15_10 <= a(15) and b(10);
        

        pp_0_11 <= a(0) and b(11);
        

        pp_1_11 <= a(1) and b(11);
        

        pp_2_11 <= a(2) and b(11);
        

        pp_3_11 <= a(3) and b(11);
        

        pp_4_11 <= a(4) and b(11);
        

        pp_5_11 <= a(5) and b(11);
        

        pp_6_11 <= a(6) and b(11);
        

        pp_7_11 <= a(7) and b(11);
        

        pp_8_11 <= a(8) and b(11);
        

        pp_9_11 <= a(9) and b(11);
        

        pp_10_11 <= a(10) and b(11);
        

        pp_11_11 <= a(11) and b(11);
        

        pp_12_11 <= a(12) and b(11);
        

        pp_13_11 <= a(13) and b(11);
        

        pp_14_11 <= a(14) and b(11);
        

        pp_15_11 <= a(15) and b(11);
        

        pp_0_12 <= a(0) and b(12);
        

        pp_1_12 <= a(1) and b(12);
        

        pp_2_12 <= a(2) and b(12);
        

        pp_3_12 <= a(3) and b(12);
        

        pp_4_12 <= a(4) and b(12);
        

        pp_5_12 <= a(5) and b(12);
        

        pp_6_12 <= a(6) and b(12);
        

        pp_7_12 <= a(7) and b(12);
        

        pp_8_12 <= a(8) and b(12);
        

        pp_9_12 <= a(9) and b(12);
        

        pp_10_12 <= a(10) and b(12);
        

        pp_11_12 <= a(11) and b(12);
        

        pp_12_12 <= a(12) and b(12);
        

        pp_13_12 <= a(13) and b(12);
        

        pp_14_12 <= a(14) and b(12);
        

        pp_15_12 <= a(15) and b(12);
        

        pp_0_13 <= a(0) and b(13);
        

        pp_1_13 <= a(1) and b(13);
        

        pp_2_13 <= a(2) and b(13);
        

        pp_3_13 <= a(3) and b(13);
        

        pp_4_13 <= a(4) and b(13);
        

        pp_5_13 <= a(5) and b(13);
        

        pp_6_13 <= a(6) and b(13);
        

        pp_7_13 <= a(7) and b(13);
        

        pp_8_13 <= a(8) and b(13);
        

        pp_9_13 <= a(9) and b(13);
        

        pp_10_13 <= a(10) and b(13);
        

        pp_11_13 <= a(11) and b(13);
        

        pp_12_13 <= a(12) and b(13);
        

        pp_13_13 <= a(13) and b(13);
        

        pp_14_13 <= a(14) and b(13);
        

        pp_15_13 <= a(15) and b(13);
        

        pp_0_14 <= a(0) and b(14);
        

        pp_1_14 <= a(1) and b(14);
        

        pp_2_14 <= a(2) and b(14);
        

        pp_3_14 <= a(3) and b(14);
        

        pp_4_14 <= a(4) and b(14);
        

        pp_5_14 <= a(5) and b(14);
        

        pp_6_14 <= a(6) and b(14);
        

        pp_7_14 <= a(7) and b(14);
        

        pp_8_14 <= a(8) and b(14);
        

        pp_9_14 <= a(9) and b(14);
        

        pp_10_14 <= a(10) and b(14);
        

        pp_11_14 <= a(11) and b(14);
        

        pp_12_14 <= a(12) and b(14);
        

        pp_13_14 <= a(13) and b(14);
        

        pp_14_14 <= a(14) and b(14);
        

        pp_15_14 <= a(15) and b(14);
        

        pp_0_15 <= a(0) and b(15);
        

        pp_1_15 <= a(1) and b(15);
        

        pp_2_15 <= a(2) and b(15);
        

        pp_3_15 <= a(3) and b(15);
        

        pp_4_15 <= a(4) and b(15);
        

        pp_5_15 <= a(5) and b(15);
        

        pp_6_15 <= a(6) and b(15);
        

        pp_7_15 <= a(7) and b(15);
        

        pp_8_15 <= a(8) and b(15);
        

        pp_9_15 <= a(9) and b(15);
        

        pp_10_15 <= a(10) and b(15);
        

        pp_11_15 <= a(11) and b(15);
        

        pp_12_15 <= a(12) and b(15);
        

        pp_13_15 <= a(13) and b(15);
        

        pp_14_15 <= a(14) and b(15);
        

        pp_15_15 <= a(15) and b(15);
        

        full_adder_1 : full_adder
            port map (
                a => pp_1_0,
                b => pp_0_1,
                Cin => '0',
                s => c(1),
                Cout => ripple_carry_1
            );
        

        full_adder_2 : full_adder
            port map (
                a => pp_2_0,
                b => sum_652062,
                Cin => ripple_carry_1,
                s => c(2),
                Cout => ripple_carry_2
            );
        

        full_adder_3 : full_adder
            port map (
                a => cout_734723,
                b => sum_454017,
                Cin => ripple_carry_2,
                s => c(3),
                Cout => ripple_carry_3
            );
        

        full_adder_4 : full_adder
            port map (
                a => cout_648852,
                b => sum_615388,
                Cin => ripple_carry_3,
                s => c(4),
                Cout => ripple_carry_4
            );
        

        full_adder_5 : full_adder
            port map (
                a => cout_622190,
                b => sum_307052,
                Cin => ripple_carry_4,
                s => c(5),
                Cout => ripple_carry_5
            );
        

        full_adder_6 : full_adder
            port map (
                a => cout_296984,
                b => sum_957721,
                Cin => ripple_carry_5,
                s => c(6),
                Cout => ripple_carry_6
            );
        

        full_adder_7 : full_adder
            port map (
                a => cout_372708,
                b => sum_910907,
                Cin => ripple_carry_6,
                s => c(7),
                Cout => ripple_carry_7
            );
        

        full_adder_8 : full_adder
            port map (
                a => cout_87182,
                b => sum_190554,
                Cin => ripple_carry_7,
                s => c(8),
                Cout => ripple_carry_8
            );
        

        full_adder_9 : full_adder
            port map (
                a => cout_901791,
                b => sum_108552,
                Cin => ripple_carry_8,
                s => c(9),
                Cout => ripple_carry_9
            );
        

        full_adder_10 : full_adder
            port map (
                a => cout_938354,
                b => sum_871398,
                Cin => ripple_carry_9,
                s => c(10),
                Cout => ripple_carry_10
            );
        

        full_adder_11 : full_adder
            port map (
                a => cout_899840,
                b => sum_748543,
                Cin => ripple_carry_10,
                s => c(11),
                Cout => ripple_carry_11
            );
        

        full_adder_12 : full_adder
            port map (
                a => cout_473235,
                b => sum_620884,
                Cin => ripple_carry_11,
                s => c(12),
                Cout => ripple_carry_12
            );
        

        full_adder_13 : full_adder
            port map (
                a => cout_502572,
                b => sum_835826,
                Cin => ripple_carry_12,
                s => c(13),
                Cout => ripple_carry_13
            );
        

        full_adder_14 : full_adder
            port map (
                a => cout_615799,
                b => sum_747437,
                Cin => ripple_carry_13,
                s => c(14),
                Cout => ripple_carry_14
            );
        

        full_adder_15 : full_adder
            port map (
                a => cout_907232,
                b => sum_408519,
                Cin => ripple_carry_14,
                s => c(15),
                Cout => ripple_carry_15
            );
        

        full_adder_16 : full_adder
            port map (
                a => cout_273843,
                b => sum_825709,
                Cin => ripple_carry_15,
                s => c(16),
                Cout => ripple_carry_16
            );
        

        full_adder_17 : full_adder
            port map (
                a => cout_593623,
                b => sum_751602,
                Cin => ripple_carry_16,
                s => c(17),
                Cout => ripple_carry_17
            );
        

        full_adder_18 : full_adder
            port map (
                a => cout_860894,
                b => sum_739794,
                Cin => ripple_carry_17,
                s => c(18),
                Cout => ripple_carry_18
            );
        

        full_adder_19 : full_adder
            port map (
                a => cout_336777,
                b => sum_422751,
                Cin => ripple_carry_18,
                s => c(19),
                Cout => ripple_carry_19
            );
        

        full_adder_20 : full_adder
            port map (
                a => cout_174675,
                b => sum_573526,
                Cin => ripple_carry_19,
                s => c(20),
                Cout => ripple_carry_20
            );
        

        full_adder_21 : full_adder
            port map (
                a => cout_622573,
                b => sum_334672,
                Cin => ripple_carry_20,
                s => c(21),
                Cout => ripple_carry_21
            );
        

        full_adder_22 : full_adder
            port map (
                a => cout_614796,
                b => sum_445479,
                Cin => ripple_carry_21,
                s => c(22),
                Cout => ripple_carry_22
            );
        

        full_adder_23 : full_adder
            port map (
                a => cout_694665,
                b => sum_873056,
                Cin => ripple_carry_22,
                s => c(23),
                Cout => ripple_carry_23
            );
        

        full_adder_24 : full_adder
            port map (
                a => cout_34362,
                b => sum_860833,
                Cin => ripple_carry_23,
                s => c(24),
                Cout => ripple_carry_24
            );
        

        full_adder_25 : full_adder
            port map (
                a => cout_288058,
                b => sum_906512,
                Cin => ripple_carry_24,
                s => c(25),
                Cout => ripple_carry_25
            );
        

        full_adder_26 : full_adder
            port map (
                a => cout_430498,
                b => sum_319921,
                Cin => ripple_carry_25,
                s => c(26),
                Cout => ripple_carry_26
            );
        

        full_adder_27 : full_adder
            port map (
                a => cout_310125,
                b => sum_777791,
                Cin => ripple_carry_26,
                s => c(27),
                Cout => ripple_carry_27
            );
        

        full_adder_28 : full_adder
            port map (
                a => cout_278529,
                b => sum_134521,
                Cin => ripple_carry_27,
                s => c(28),
                Cout => ripple_carry_28
            );
        

        full_adder_29 : full_adder
            port map (
                a => cout_907380,
                b => sum_453295,
                Cin => ripple_carry_28,
                s => c(29),
                Cout => ripple_carry_29
            );
        

        full_adder_30 : full_adder
            port map (
                a => pp_15_15,
                b => cout_505573,
                Cin => ripple_carry_29,
                s => c(30),
                Cout => ripple_carry_30
            );
        
c(0) <= pp_0_0;

end Behavioral;
